// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION

`include "jpc_global.v"

`define	MAX_PATH			256
module tb();

	parameter  FRAME_WIDTH = 112;
	parameter  FRAME_HEIGHT = 48;
	parameter  SIM_FRAMES = 2;
	reg						rstn;
	reg						clk;
	reg						ee_clk;
	
	wire		rstn_ee = rstn;
	initial begin
		rstn = `RESET_ACTIVE;
		#(`RESET_DELAY); 
		$display("T%d rstn done#############################", $time);
		rstn = `RESET_IDLE;
	end
	
	initial begin
		clk = 1;
		forever begin
			clk = ~clk;
			#(`CLK_PERIOD_DIV2);
		end
	end
	
	initial begin
		ee_clk = 1;
		forever begin
			ee_clk = ~ee_clk;
			#(`EE_CLOCK_PERIOD_DIV2);
		end
	end
	
	reg		gt_ref_clk;
	initial begin
		gt_ref_clk = 1;
		forever begin
			gt_ref_clk = ~gt_ref_clk;
			#(`GT_REF_CLOCK_PERIOD_DIV2);
		end
	end
	
	reg			[15:0]			frame_width_0;
	reg			[15:0]			frame_height_0;
	reg			[31:0]			pic_to_sim;
	reg		[`MAX_PATH*8-1:0]	sequence_name_0;

	itf itf(clk);

	wire					go = itf.go;
	initial begin
		itf.init();
		#(`RESET_DELAY)
		#(`RESET_DELAY)
		// itf.start();
		itf.drive();
		//itf.drive_a_frame();
	end	




	wire	[13:0]			aa_src_rom;
	wire	[`W2:0]			qa_src_rom;

	
	src_rom src_rom(
		.clk			(clk),
		.rstn			(rstn),
		.aa				(aa_src_rom),
		.cena			(cena_src_rom),
		.qa				(qa_src_rom)
		);
		
		

	wire	[15:0]	num_tile_in_pic = 16;
	wire	[15:0]	pic_width = `TILE_WIDTH * 4;
	wire	[15:0]	pic_height = `TILE_WIDTH * 4;
	wire	[ 3:0]	ndecomp = 1;

	
	wire	 				data_valid;
	wire	[7:0]			data_out;
	
	reg					doing_enc;
	reg		[15:0]		tile_cnt;
	wire				enc_go;
	
	wire		unset_doing_enc = enc_go & tile_cnt==num_tile_in_pic-1;
	
	always @(`CLK_RST_EDGE)
		if (`RST)			tile_cnt <= 0;
		else if (go)		tile_cnt <= 0;
		else if (enc_go)	tile_cnt <= tile_cnt + 1;

	wire	first_tile_f = tile_cnt ==0;
	wire	last_tile_f = tile_cnt==num_tile_in_pic-1;
	
	always @(`CLK_RST_EDGE)
		if (`RST)					doing_enc <= 0;
		else if (go)				doing_enc <= 1;
		else if (unset_doing_enc)	doing_enc <= 0;
	
	wire	enc_busy;
	assign	enc_go = doing_enc & !enc_busy;

	jpc_core jpc_core(
		.clk			(clk),
		.rstn			(rstn),

		.go				(enc_go),
		.first_tile_f	(first_tile_f),
		.last_tile_f	(last_tile_f),
		
		.pic_width		(pic_width),
		.pic_height		(pic_height),
		.ndecomp		(ndecomp),

		.cena_src_buf	(cena_src_rom),
		.aa_src_buf		(aa_src_rom),
		.qa_src_buf		(qa_src_rom),


		.byte_out_f		(data_valid),
		.byte_out		(data_out),

		.busy			(enc_busy),
		.pic_ready		(pic_ready),
		.ready			()
		);

	always @(`CLK_EDGE)
		if (pic_ready) begin
			$display("======= encode pic done =========");
			#200 $finish();
		end

	`DELAYEN8(data_out, 7, data_valid)
	reg		[15:0]	pic_data_cnt;
	always @(`CLK_RST_EDGE)
		if (`RST)					pic_data_cnt <= 0;
		else if (data_valid)		pic_data_cnt <= pic_data_cnt +1;
	wire 	[31:0]	pic_words = { data_out, 
									data_out_d1, 
									data_out_d2, 
									data_out_d3
								};
	reg		[`MAX_PATH*8-1:0]	pic_dsc = "enc.jpc";
	integer						fds_pic_dsc;
	initial
		fds_pic_dsc = $fopen(pic_dsc, "wb");
	always @(`CLK_RST_EDGE)
		if (data_valid && pic_data_cnt[1:0]==2'b11) begin
			$fwrite(fds_pic_dsc, "%u", pic_words);
		end							

`ifdef DUMP_FSDB 
	initial begin
	$fsdbDumpfile("fsdb/xx.fsdb");
	//$fsdbDumpvars();
	$fsdbDumpvars(5, tb);
	end
`endif
	
endmodule




module src_rom(
	input			clk,
	input			rstn,
	input	[13:0]	aa,
	input			cena,
	output reg		[`W2:0]	qa
	);
	logic [0:`TILE_WIDTH*`TILE_WIDTH-1][31:0] mem	 = {
 -66, 	 -70, 	 -74, 	 -80, 	 -76, 	 -51, 	 -43, 	 -39, 	 -38, 	 -37, 	 -36, 	 -29, 	 -60, 	 -67, 	 -64, 	 -59, 	 -47, 	 -22, 	  30, 	  34, 	  38, 	  35, 	  35, 	  34, 	  33, 	  32, 	  32, 	  31, 	  27, 	  -7, 	 -76, 	 -81, 	 -82, 	 -86, 	 -85, 	 -86, 	 -84, 	 -84, 	 -84, 	 -82, 	 -76, 	 -75, 	 -73, 	 -74, 	 -74, 	 -72, 	 -70, 	 -68, 	 -67, 	 -65, 	 -63, 	 -60, 	 -58, 	 -58, 	 -56, 	 -56, 	 -52, 	 -55, 	 -60, 	 -61, 	 -58, 	 -57, 	 -57, 	 -57, 		 -53, 	 -66, 	 -50, 	 -52, 	 -67, 	 -71, 	 -70, 	 -70, 	 -70, 	 -73, 	 -67, 	 -46, 	 -71, 	 -83, 	 -83, 	 -82, 	 -65, 	 -49, 	 -31, 	 -74, 	 -85, 	 -85, 	 -87, 	 -86, 	 -86, 	 -86, 	 -86, 	 -84, 	 -85, 	 -86, 	 -86, 	 -85, 	 -85, 	 -85, 	 -84, 	 -86, 	 -86, 	 -87, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -87, 	 -85, 	 -85, 	 -85, 	 -80, 	 -77, 	 -80, 	 -82, 	 -80, 	 -77, 	 -74, 	 -73, 	 -75, 	 -73, 	 -71, 	 -72, 	 -72, 	
 -66, 	 -70, 	 -75, 	 -77, 	 -77, 	 -52, 	 -40, 	 -37, 	 -35, 	 -41, 	 -30, 	 -30, 	 -59, 	 -67, 	 -64, 	 -55, 	 -46, 	 -23, 	  27, 	  33, 	  38, 	  35, 	  35, 	  37, 	  36, 	  38, 	  36, 	  34, 	  32, 	  -6, 	 -77, 	 -82, 	 -82, 	 -83, 	 -83, 	 -86, 	 -84, 	 -84, 	 -83, 	 -83, 	 -77, 	 -75, 	 -73, 	 -75, 	 -74, 	 -72, 	 -69, 	 -68, 	 -67, 	 -63, 	 -62, 	 -60, 	 -60, 	 -56, 	 -54, 	 -54, 	 -53, 	 -58, 	 -63, 	 -57, 	 -57, 	 -54, 	 -60, 	 -58, 		 -69, 	 -78, 	 -79, 	 -65, 	 -64, 	 -72, 	 -74, 	 -74, 	 -71, 	 -71, 	 -68, 	 -48, 	 -55, 	 -84, 	 -83, 	 -86, 	 -81, 	 -64, 	 -42, 	 -64, 	 -84, 	 -88, 	 -88, 	 -86, 	 -86, 	 -86, 	 -85, 	 -84, 	 -87, 	 -85, 	 -85, 	 -86, 	 -85, 	 -86, 	 -87, 	 -85, 	 -86, 	 -87, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -81, 	 -85, 	 -85, 	 -81, 	 -75, 	 -73, 	 -82, 	 -80, 	 -76, 	 -71, 	 -68, 	 -65, 	 -64, 	 -66, 	 -69, 	 -72, 	
 -75, 	 -74, 	 -76, 	 -79, 	 -77, 	 -48, 	 -39, 	 -37, 	 -39, 	 -37, 	 -35, 	 -29, 	 -61, 	 -61, 	 -57, 	 -59, 	 -54, 	 -46, 	  -8, 	  14, 	  19, 	  21, 	  26, 	  31, 	  32, 	  35, 	  34, 	  35, 	  29, 	  -6, 	 -75, 	 -81, 	 -78, 	 -86, 	 -83, 	 -84, 	 -86, 	 -84, 	 -82, 	 -80, 	 -75, 	 -74, 	 -75, 	 -73, 	 -71, 	 -74, 	 -69, 	 -71, 	 -67, 	 -66, 	 -63, 	 -61, 	 -59, 	 -54, 	 -56, 	 -56, 	 -55, 	 -61, 	 -63, 	 -61, 	 -58, 	 -59, 	 -59, 	 -60, 		 -64, 	 -72, 	 -77, 	 -65, 	 -70, 	 -74, 	 -79, 	 -76, 	 -71, 	 -62, 	 -53, 	 -48, 	 -49, 	 -64, 	 -78, 	 -82, 	 -85, 	 -79, 	 -61, 	 -52, 	 -78, 	 -87, 	 -86, 	 -83, 	 -85, 	 -87, 	 -85, 	 -86, 	 -86, 	 -85, 	 -85, 	 -86, 	 -85, 	 -85, 	 -85, 	 -86, 	 -87, 	 -87, 	 -85, 	 -86, 	 -86, 	 -86, 	 -86, 	 -87, 	 -87, 	 -85, 	 -86, 	 -85, 	 -80, 	 -80, 	 -82, 	 -82, 	 -76, 	 -69, 	 -73, 	 -72, 	 -66, 	 -52, 	  -8, 	  -1, 	   1, 	  -9, 	 -47, 	 -69, 	
 -82, 	 -80, 	 -76, 	 -80, 	 -76, 	 -48, 	 -36, 	 -37, 	 -35, 	 -36, 	 -34, 	 -23, 	 -54, 	 -69, 	 -67, 	 -70, 	 -69, 	 -67, 	 -61, 	 -53, 	 -44, 	 -37, 	 -35, 	 -26, 	 -25, 	 -17, 	  -6, 	   4, 	  14, 	  -4, 	 -32, 	 -39, 	 -49, 	 -60, 	 -66, 	 -74, 	 -76, 	 -79, 	 -82, 	 -80, 	 -79, 	 -73, 	 -72, 	 -71, 	 -71, 	 -70, 	 -70, 	 -69, 	 -66, 	 -66, 	 -63, 	 -59, 	 -56, 	 -56, 	 -52, 	 -54, 	 -57, 	 -65, 	 -65, 	 -56, 	 -57, 	 -56, 	 -60, 	 -63, 		 -63, 	 -57, 	 -53, 	 -51, 	 -59, 	 -60, 	 -65, 	 -57, 	 -38, 	 -28, 	 -22, 	 -44, 	 -37, 	 -34, 	 -66, 	 -83, 	 -83, 	 -86, 	 -79, 	 -56, 	 -62, 	 -75, 	 -86, 	 -86, 	 -86, 	 -86, 	 -85, 	 -84, 	 -85, 	 -85, 	 -85, 	 -86, 	 -85, 	 -85, 	 -85, 	 -86, 	 -87, 	 -87, 	 -85, 	 -86, 	 -86, 	 -86, 	 -86, 	 -87, 	 -87, 	 -85, 	 -86, 	 -85, 	 -76, 	 -81, 	 -82, 	 -82, 	 -81, 	 -78, 	 -72, 	 -56, 	 -51, 	 -52, 	 -41, 	 -42, 	 -63, 	 -70, 	 -70, 	 -70, 	
 -85, 	 -80, 	 -77, 	 -77, 	 -75, 	 -45, 	 -36, 	 -36, 	 -38, 	 -34, 	 -32, 	 -31, 	 -44, 	 -62, 	 -64, 	 -65, 	 -67, 	 -70, 	 -71, 	 -72, 	 -74, 	 -72, 	 -72, 	 -69, 	 -63, 	 -60, 	 -57, 	 -50, 	 -45, 	 -35, 	 -33, 	 -27, 	 -27, 	 -25, 	 -25, 	 -29, 	 -28, 	 -34, 	 -37, 	 -38, 	 -42, 	 -39, 	 -38, 	 -46, 	 -48, 	 -54, 	 -60, 	 -64, 	 -65, 	 -64, 	 -59, 	 -61, 	 -61, 	 -53, 	 -53, 	 -53, 	 -55, 	 -67, 	 -64, 	 -58, 	 -57, 	 -58, 	 -59, 	 -60, 		 -61, 	 -56, 	 -44, 	 -42, 	 -50, 	 -37, 	 -31, 	 -17, 	   6, 	 -16, 	 -17, 	 -43, 	 -35, 	 -24, 	 -36, 	 -72, 	 -80, 	 -85, 	 -84, 	 -76, 	 -58, 	 -65, 	 -86, 	 -84, 	 -84, 	 -86, 	 -85, 	 -85, 	 -84, 	 -85, 	 -85, 	 -85, 	 -85, 	 -86, 	 -85, 	 -86, 	 -87, 	 -87, 	 -85, 	 -86, 	 -86, 	 -86, 	 -86, 	 -87, 	 -87, 	 -86, 	 -86, 	 -82, 	 -78, 	 -85, 	 -85, 	 -85, 	 -84, 	 -78, 	 -75, 	 -63, 	 -61, 	 -61, 	 -41, 	 -40, 	 -53, 	 -79, 	 -80, 	 -78, 	
 -83, 	 -76, 	 -73, 	 -72, 	 -65, 	 -36, 	 -37, 	 -31, 	 -34, 	 -31, 	 -32, 	 -12, 	 -11, 	 -15, 	 -26, 	 -39, 	 -50, 	 -53, 	 -62, 	 -64, 	 -63, 	 -65, 	 -72, 	 -70, 	 -75, 	 -75, 	 -77, 	 -76, 	 -72, 	 -66, 	 -64, 	 -61, 	 -54, 	 -51, 	 -43, 	 -42, 	 -38, 	 -34, 	 -30, 	 -29, 	 -29, 	 -20, 	 -16, 	 -16, 	 -11, 	  -7, 	  -8, 	 -13, 	 -18, 	 -29, 	 -45, 	 -51, 	 -52, 	 -49, 	 -52, 	 -52, 	 -54, 	 -65, 	 -62, 	 -58, 	 -57, 	 -59, 	 -58, 	 -58, 		 -57, 	 -56, 	 -42, 	 -41, 	 -43, 	 -33, 	 -27, 	  -8, 	  10, 	 -11, 	 -16, 	 -43, 	 -35, 	 -20, 	 -23, 	 -44, 	 -78, 	 -84, 	 -84, 	 -84, 	 -76, 	 -63, 	 -72, 	 -83, 	 -88, 	 -84, 	 -85, 	 -86, 	 -82, 	 -79, 	 -85, 	 -85, 	 -85, 	 -86, 	 -85, 	 -87, 	 -88, 	 -87, 	 -87, 	 -86, 	 -85, 	 -85, 	 -86, 	 -85, 	 -87, 	 -86, 	 -80, 	 -79, 	 -77, 	 -85, 	 -85, 	 -86, 	 -85, 	 -77, 	 -79, 	 -78, 	 -74, 	 -74, 	 -65, 	 -66, 	 -57, 	 -65, 	 -76, 	 -74, 	
 -72, 	 -73, 	 -69, 	 -62, 	 -46, 	 -32, 	 -29, 	 -28, 	 -29, 	 -29, 	 -28, 	 -32, 	 -31, 	 -31, 	 -28, 	 -24, 	 -22, 	 -15, 	  -9, 	  -9, 	 -17, 	 -33, 	 -40, 	 -54, 	 -59, 	 -64, 	 -65, 	 -70, 	 -70, 	 -77, 	 -75, 	 -75, 	 -78, 	 -70, 	 -68, 	 -63, 	 -62, 	 -56, 	 -54, 	 -49, 	 -42, 	 -26, 	 -25, 	 -23, 	 -16, 	  -8, 	  -7, 	  -4, 	  -5, 	  -3, 	   0, 	   3, 	   0, 	 -14, 	 -26, 	 -40, 	 -48, 	 -61, 	 -58, 	 -56, 	 -57, 	 -59, 	 -59, 	 -57, 		 -59, 	 -49, 	 -38, 	 -45, 	 -43, 	 -27, 	 -25, 	  -7, 	   8, 	 -14, 	 -19, 	 -42, 	 -32, 	 -18, 	 -18, 	 -24, 	 -48, 	 -79, 	 -79, 	 -83, 	 -85, 	 -75, 	 -59, 	 -76, 	 -86, 	 -85, 	 -84, 	 -84, 	 -77, 	 -68, 	 -82, 	 -85, 	 -84, 	 -85, 	 -88, 	 -85, 	 -87, 	 -81, 	 -85, 	 -85, 	 -86, 	 -84, 	 -85, 	 -85, 	 -85, 	 -87, 	 -84, 	 -81, 	 -84, 	 -85, 	 -85, 	 -85, 	 -81, 	 -79, 	 -77, 	 -76, 	 -80, 	 -78, 	 -74, 	 -82, 	 -82, 	 -79, 	 -80, 	 -75, 	
 -69, 	 -60, 	 -34, 	 -18, 	  -6, 	   1, 	   0, 	   2, 	   6, 	  12, 	   4, 	  -6, 	 -18, 	 -28, 	 -31, 	 -35, 	 -29, 	 -34, 	 -33, 	 -34, 	 -33, 	 -32, 	 -27, 	 -20, 	 -13, 	 -16, 	 -17, 	 -25, 	 -35, 	 -48, 	 -60, 	 -66, 	 -67, 	 -68, 	 -73, 	 -72, 	 -75, 	 -71, 	 -71, 	 -67, 	 -61, 	 -47, 	 -39, 	 -34, 	 -32, 	 -26, 	 -23, 	 -14, 	 -14, 	 -14, 	  -8, 	   5, 	   6, 	   5, 	  14, 	  11, 	   5, 	  -6, 	 -26, 	 -38, 	 -47, 	 -52, 	 -49, 	 -52, 		 -50, 	 -41, 	 -44, 	 -43, 	 -38, 	 -26, 	 -21, 	  -5, 	   4, 	 -45, 	 -40, 	 -40, 	 -34, 	 -17, 	 -19, 	 -21, 	 -24, 	 -56, 	 -80, 	 -81, 	 -83, 	 -81, 	 -75, 	 -58, 	 -76, 	 -82, 	 -83, 	 -82, 	 -81, 	 -69, 	 -78, 	 -86, 	 -85, 	 -84, 	 -83, 	 -86, 	 -84, 	 -83, 	 -82, 	 -84, 	 -86, 	 -84, 	 -85, 	 -85, 	 -85, 	 -86, 	 -86, 	 -83, 	 -84, 	 -85, 	 -85, 	 -85, 	 -83, 	 -82, 	 -80, 	 -76, 	 -74, 	 -79, 	 -82, 	 -81, 	 -81, 	 -77, 	 -74, 	 -71, 	
 -14, 	   7, 	  33, 	  36, 	  37, 	  34, 	  35, 	  30, 	  47, 	  46, 	  31, 	  20, 	   3, 	 -17, 	 -30, 	 -28, 	 -26, 	 -26, 	 -29, 	 -31, 	 -34, 	 -32, 	 -33, 	 -31, 	 -32, 	 -28, 	 -34, 	 -30, 	 -27, 	 -24, 	 -20, 	 -19, 	 -21, 	 -26, 	 -34, 	 -49, 	 -58, 	 -63, 	 -66, 	 -65, 	 -65, 	 -57, 	 -57, 	 -51, 	 -46, 	 -41, 	 -32, 	 -24, 	 -20, 	 -10, 	  -5, 	  -1, 	   3, 	   5, 	   5, 	   1, 	   2, 	   1, 	   2, 	  -2, 	  -8, 	 -20, 	 -14, 	 -21, 		 -17, 	 -19, 	 -23, 	 -18, 	 -20, 	 -27, 	 -22, 	  -4, 	   6, 	 -50, 	 -51, 	 -37, 	 -34, 	 -16, 	 -16, 	 -21, 	 -23, 	 -31, 	 -63, 	 -78, 	 -82, 	 -85, 	 -80, 	 -71, 	 -61, 	 -74, 	 -82, 	 -83, 	 -81, 	 -56, 	 -73, 	 -88, 	 -83, 	 -86, 	 -82, 	 -84, 	 -86, 	 -80, 	 -82, 	 -84, 	 -86, 	 -84, 	 -85, 	 -87, 	 -86, 	 -85, 	 -85, 	 -85, 	 -79, 	 -77, 	 -70, 	 -78, 	 -82, 	 -80, 	 -82, 	 -79, 	 -78, 	 -80, 	 -77, 	 -78, 	 -75, 	 -72, 	 -69, 	 -71, 	
  47, 	  52, 	  60, 	  62, 	  61, 	  63, 	  63, 	  46, 	  44, 	  53, 	  42, 	  39, 	  25, 	  11, 	 -13, 	 -27, 	 -29, 	 -33, 	 -42, 	 -40, 	 -39, 	 -35, 	 -33, 	 -27, 	 -26, 	 -26, 	 -28, 	 -31, 	 -30, 	 -30, 	 -30, 	 -30, 	 -29, 	 -29, 	 -24, 	 -20, 	 -19, 	 -14, 	 -18, 	 -29, 	 -37, 	 -47, 	 -51, 	 -56, 	 -52, 	 -40, 	 -34, 	 -21, 	 -16, 	 -17, 	 -10, 	 -12, 	  -6, 	 -11, 	  -8, 	 -11, 	 -15, 	 -23, 	 -24, 	 -25, 	 -27, 	 -29, 	 -33, 	 -35, 		 -30, 	 -32, 	 -35, 	 -31, 	 -27, 	 -15, 	 -24, 	  -5, 	   9, 	 -12, 	 -32, 	 -39, 	 -28, 	 -18, 	 -19, 	 -18, 	 -19, 	 -22, 	 -34, 	 -73, 	 -78, 	 -81, 	 -85, 	 -78, 	 -70, 	 -60, 	 -65, 	 -77, 	 -77, 	 -55, 	 -53, 	 -82, 	 -83, 	 -80, 	 -84, 	 -83, 	 -85, 	 -79, 	 -84, 	 -84, 	 -83, 	 -83, 	 -85, 	 -84, 	 -83, 	 -83, 	 -84, 	 -81, 	 -72, 	 -73, 	 -69, 	 -69, 	 -74, 	 -75, 	 -75, 	 -78, 	 -81, 	 -79, 	 -80, 	 -81, 	 -78, 	 -73, 	 -76, 	 -71, 	
  59, 	  59, 	  65, 	  67, 	  67, 	  67, 	  67, 	  66, 	  63, 	  60, 	  61, 	  55, 	  52, 	  46, 	  47, 	  37, 	  30, 	  18, 	   5, 	 -10, 	 -20, 	 -23, 	 -31, 	 -33, 	 -41, 	 -42, 	 -36, 	 -33, 	 -30, 	 -22, 	 -24, 	 -26, 	 -25, 	 -31, 	 -26, 	 -31, 	 -28, 	 -31, 	 -27, 	 -26, 	 -19, 	 -12, 	  -3, 	  -3, 	  -8, 	  -9, 	 -20, 	 -30, 	 -35, 	 -38, 	 -38, 	 -31, 	 -23, 	 -14, 	 -16, 	 -14, 	 -24, 	 -24, 	 -26, 	 -26, 	 -25, 	 -25, 	 -26, 	 -26, 		 -28, 	 -26, 	 -25, 	 -25, 	 -18, 	  -9, 	  -9, 	   0, 	  12, 	  -5, 	 -27, 	 -34, 	 -29, 	 -15, 	 -16, 	 -19, 	 -22, 	 -18, 	 -24, 	 -36, 	 -75, 	 -80, 	 -81, 	 -85, 	 -81, 	 -73, 	 -62, 	 -70, 	 -74, 	 -57, 	 -57, 	 -78, 	 -81, 	 -81, 	 -81, 	 -82, 	 -79, 	 -84, 	 -81, 	 -83, 	 -83, 	 -83, 	 -82, 	 -83, 	 -82, 	 -81, 	 -81, 	 -82, 	 -69, 	 -66, 	 -60, 	 -55, 	 -59, 	 -63, 	 -67, 	 -74, 	 -78, 	 -79, 	 -70, 	 -62, 	 -66, 	 -69, 	 -69, 	 -69, 	
  58, 	  61, 	  59, 	  62, 	  61, 	  63, 	  64, 	  67, 	  65, 	  65, 	  66, 	  68, 	  67, 	  61, 	  65, 	  61, 	  60, 	  56, 	  50, 	  49, 	  44, 	  46, 	  40, 	  27, 	  18, 	   3, 	  -7, 	 -21, 	 -28, 	 -35, 	 -41, 	 -41, 	 -44, 	 -38, 	 -32, 	 -26, 	 -24, 	 -25, 	 -27, 	 -26, 	 -26, 	 -22, 	 -19, 	 -16, 	 -12, 	  -6, 	  -4, 	   4, 	  13, 	  14, 	  17, 	  24, 	  32, 	  46, 	  69, 	  18, 	   9, 	   7, 	  11, 	  13, 	   5, 	   4, 	  -3, 	  -6, 		 -13, 	 -20, 	 -18, 	 -22, 	 -23, 	 -20, 	  -5, 	  17, 	  15, 	  -5, 	 -25, 	 -31, 	 -20, 	 -15, 	 -17, 	 -15, 	 -16, 	 -19, 	 -20, 	 -26, 	 -47, 	 -76, 	 -79, 	 -82, 	 -86, 	 -78, 	 -73, 	 -63, 	 -71, 	 -51, 	 -48, 	 -76, 	 -78, 	 -78, 	 -81, 	 -79, 	 -80, 	 -76, 	 -76, 	 -74, 	 -71, 	 -66, 	 -64, 	 -62, 	 -57, 	 -54, 	 -53, 	 -45, 	 -39, 	 -35, 	 -33, 	 -19, 	 -23, 	 -27, 	 -35, 	 -34, 	 -36, 	 -34, 	 -39, 	 -36, 	 -35, 	 -41, 	 -40, 	 -31, 	
  48, 	  47, 	  49, 	  51, 	  53, 	  52, 	  58, 	  61, 	  59, 	  59, 	  62, 	  62, 	  63, 	  63, 	  64, 	  65, 	  62, 	  62, 	  62, 	  61, 	  60, 	  63, 	  60, 	  58, 	  57, 	  57, 	  50, 	  46, 	  40, 	  34, 	  18, 	   4, 	 -12, 	 -25, 	 -33, 	 -35, 	 -40, 	 -39, 	 -37, 	 -30, 	 -21, 	  -9, 	  -8, 	  -7, 	  -7, 	  -6, 	  -8, 	  -6, 	  -4, 	  -2, 	  -2, 	   0, 	   0, 	   4, 	  14, 	   0, 	   1, 	  -2, 	   0, 	   0, 	  -1, 	   1, 	   1, 	   4, 		   5, 	   5, 	  11, 	  12, 	  10, 	   7, 	  17, 	  20, 	   4, 	   2, 	 -24, 	 -26, 	 -20, 	 -20, 	 -25, 	 -24, 	 -30, 	 -33, 	 -37, 	 -39, 	 -47, 	 -67, 	 -77, 	 -77, 	 -80, 	 -84, 	 -78, 	 -70, 	 -50, 	 -22, 	 -15, 	 -32, 	 -35, 	 -32, 	 -32, 	 -33, 	 -29, 	 -24, 	 -25, 	 -25, 	 -25, 	 -25, 	 -27, 	 -28, 	 -31, 	 -35, 	 -37, 	 -35, 	 -34, 	 -33, 	 -32, 	 -30, 	 -28, 	 -32, 	 -31, 	 -38, 	 -42, 	 -38, 	 -36, 	 -34, 	 -33, 	 -33, 	 -36, 	 -37, 	
  39, 	  39, 	  42, 	  40, 	  39, 	  47, 	  44, 	  47, 	  49, 	  51, 	  53, 	  56, 	  57, 	  56, 	  59, 	  57, 	  57, 	  56, 	  56, 	  58, 	  58, 	  58, 	  55, 	  55, 	  55, 	  55, 	  52, 	  52, 	  48, 	  46, 	  49, 	  45, 	  44, 	  46, 	  43, 	  34, 	  18, 	   7, 	 -13, 	 -21, 	 -10, 	   2, 	   3, 	   5, 	   7, 	  12, 	  13, 	  14, 	  18, 	  15, 	  16, 	  17, 	  13, 	  11, 	  10, 	   9, 	   5, 	  -3, 	  -2, 	  -2, 	  -4, 	  -8, 	  -6, 	  -7, 		  -7, 	  -7, 	  -9, 	  -9, 	  -5, 	  -5, 	  -5, 	  -3, 	   0, 	  -3, 	 -27, 	 -27, 	 -13, 	  -6, 	  -4, 	 -10, 	 -14, 	 -15, 	 -10, 	 -10, 	 -10, 	 -26, 	 -67, 	 -79, 	 -83, 	 -80, 	 -81, 	 -75, 	 -67, 	 -44, 	 -38, 	 -42, 	 -38, 	 -38, 	 -43, 	 -46, 	 -46, 	 -47, 	 -52, 	 -52, 	 -53, 	 -54, 	 -58, 	 -60, 	 -63, 	 -65, 	 -66, 	 -65, 	 -65, 	 -66, 	 -62, 	 -61, 	 -59, 	 -64, 	 -68, 	 -72, 	 -77, 	 -77, 	 -77, 	 -77, 	 -75, 	 -76, 	 -76, 	 -78, 	
  30, 	  31, 	  29, 	  33, 	  37, 	  41, 	  43, 	  47, 	  46, 	  42, 	  42, 	  41, 	  45, 	  45, 	  50, 	  51, 	  54, 	  55, 	  54, 	  55, 	  55, 	  58, 	  54, 	  54, 	  55, 	  54, 	  55, 	  52, 	  51, 	  49, 	  51, 	  48, 	  51, 	  50, 	  49, 	  41, 	  47, 	  44, 	  46, 	  48, 	  53, 	  58, 	  57, 	  53, 	  52, 	  50, 	  46, 	  41, 	  40, 	  32, 	  33, 	  31, 	  25, 	  21, 	  24, 	  25, 	  20, 	  14, 	  14, 	  11, 	   5, 	   5, 	   8, 	   7, 		   9, 	   9, 	   5, 	   6, 	   6, 	   3, 	   0, 	   9, 	  -1, 	 -11, 	 -27, 	 -26, 	  -2, 	  37, 	  24, 	  10, 	   9, 	  -6, 	 -14, 	 -32, 	 -33, 	 -27, 	 -40, 	 -67, 	 -81, 	 -81, 	 -82, 	 -80, 	 -78, 	 -70, 	 -66, 	 -65, 	 -66, 	 -68, 	 -63, 	 -69, 	 -65, 	 -63, 	 -66, 	 -66, 	 -70, 	 -69, 	 -67, 	 -69, 	 -68, 	 -70, 	 -72, 	 -71, 	 -73, 	 -76, 	 -72, 	 -76, 	 -78, 	 -77, 	 -80, 	 -78, 	 -81, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -84, 	 -83, 	
  30, 	  30, 	  26, 	  26, 	  30, 	  28, 	  33, 	  35, 	  40, 	  42, 	  44, 	  47, 	  50, 	  50, 	  51, 	  50, 	  48, 	  51, 	  53, 	  60, 	  58, 	  60, 	  57, 	  58, 	  58, 	  59, 	  58, 	  58, 	  59, 	  57, 	  57, 	  57, 	  60, 	  58, 	  59, 	  58, 	  53, 	  54, 	  49, 	  48, 	  50, 	  54, 	  55, 	  57, 	  61, 	  56, 	  59, 	  61, 	  60, 	  63, 	  60, 	  61, 	  63, 	  60, 	  57, 	  56, 	  54, 	  50, 	  48, 	  46, 	  36, 	  30, 	  27, 	  23, 		  22, 	  17, 	  17, 	  18, 	  18, 	  25, 	  19, 	   7, 	  -5, 	  -7, 	  -8, 	 -28, 	   1, 	  32, 	  38, 	  28, 	  31, 	  19, 	   8, 	  13, 	   9, 	  14, 	   6, 	  -9, 	 -43, 	 -61, 	 -73, 	 -79, 	 -75, 	 -81, 	 -75, 	 -79, 	 -78, 	 -77, 	 -76, 	 -74, 	 -78, 	 -75, 	 -70, 	 -68, 	 -68, 	 -65, 	 -59, 	 -57, 	 -51, 	 -47, 	 -44, 	 -61, 	 -75, 	 -76, 	 -76, 	 -76, 	 -73, 	 -77, 	 -74, 	 -73, 	 -76, 	 -74, 	 -76, 	 -75, 	 -78, 	 -78, 	 -76, 	 -76, 	
  32, 	  29, 	  34, 	  26, 	  26, 	  28, 	  31, 	  25, 	  28, 	  28, 	  25, 	  26, 	  35, 	  39, 	  44, 	  46, 	  48, 	  54, 	  53, 	  51, 	  53, 	  54, 	  53, 	  62, 	  58, 	  61, 	  63, 	  62, 	  63, 	  62, 	  57, 	  62, 	  63, 	  63, 	  60, 	  64, 	  62, 	  63, 	  64, 	  59, 	  59, 	  60, 	  61, 	  60, 	  63, 	  61, 	  58, 	  60, 	  59, 	  60, 	  58, 	  58, 	  55, 	  57, 	  58, 	  55, 	  56, 	  56, 	  55, 	  54, 	  52, 	  53, 	  53, 	  51, 		  49, 	  48, 	  49, 	  49, 	  50, 	  53, 	  45, 	  32, 	  10, 	   3, 	 -15, 	 -47, 	 -12, 	  44, 	  39, 	  34, 	  32, 	  22, 	  23, 	  21, 	  20, 	  17, 	  12, 	   6, 	  -1, 	  -7, 	 -17, 	 -39, 	 -64, 	 -69, 	 -71, 	 -73, 	 -74, 	 -73, 	 -73, 	 -76, 	 -72, 	 -49, 	  -7, 	  -7, 	  -3, 	   0, 	   3, 	   4, 	   7, 	  11, 	  13, 	   3, 	 -39, 	 -61, 	 -63, 	 -65, 	 -61, 	 -56, 	 -55, 	 -57, 	 -60, 	 -64, 	 -66, 	 -71, 	 -69, 	 -69, 	 -69, 	 -77, 	
  23, 	  24, 	  25, 	  31, 	  26, 	  24, 	  16, 	  20, 	  23, 	  25, 	  31, 	  36, 	  31, 	  38, 	  37, 	  34, 	  31, 	  29, 	  43, 	  43, 	  44, 	  45, 	  50, 	  49, 	  53, 	  55, 	  54, 	  58, 	  51, 	  43, 	  52, 	  57, 	  63, 	  64, 	  64, 	  64, 	  66, 	  66, 	  64, 	  63, 	  64, 	  64, 	  64, 	  66, 	  63, 	  62, 	  63, 	  62, 	  63, 	  61, 	  59, 	  61, 	  60, 	  56, 	  60, 	  59, 	  60, 	  55, 	  56, 	  55, 	  54, 	  53, 	  53, 	  48, 		  53, 	  53, 	  54, 	  59, 	  59, 	  57, 	  51, 	  49, 	  25, 	  -6, 	 -23, 	 -10, 	  -2, 	   8, 	   4, 	  -6, 	  -7, 	 -17, 	 -27, 	 -21, 	 -33, 	 -35, 	 -43, 	 -45, 	 -48, 	 -46, 	 -40, 	 -50, 	 -55, 	 -60, 	 -56, 	 -61, 	 -58, 	 -61, 	 -62, 	 -58, 	 -63, 	 -71, 	 -61, 	  -8, 	   8, 	  13, 	  10, 	  12, 	  12, 	  18, 	  18, 	  17, 	   7, 	 -34, 	 -48, 	 -50, 	 -53, 	 -53, 	 -56, 	 -56, 	 -56, 	 -61, 	 -61, 	 -60, 	 -58, 	 -56, 	 -60, 	 -68, 	
  24, 	  28, 	  35, 	  32, 	  31, 	  27, 	  33, 	  33, 	  35, 	  28, 	  30, 	  33, 	  33, 	  32, 	  34, 	  32, 	  25, 	  28, 	  21, 	  20, 	  18, 	   9, 	  15, 	  26, 	  22, 	  31, 	  35, 	  33, 	  33, 	  34, 	  37, 	  42, 	  44, 	  49, 	  58, 	  57, 	  60, 	  65, 	  68, 	  69, 	  69, 	  64, 	  62, 	  62, 	  65, 	  67, 	  65, 	  67, 	  63, 	  63, 	  61, 	  64, 	  67, 	  67, 	  66, 	  67, 	  66, 	  66, 	  64, 	  62, 	  64, 	  64, 	  62, 	  61, 		  57, 	  58, 	  57, 	  59, 	  61, 	  61, 	  61, 	  60, 	  51, 	  53, 	  47, 	  35, 	  20, 	  -3, 	 -29, 	 -42, 	 -44, 	 -53, 	 -48, 	 -53, 	 -50, 	 -52, 	 -51, 	 -51, 	 -43, 	 -39, 	 -45, 	 -55, 	 -54, 	 -57, 	 -56, 	 -57, 	 -56, 	 -53, 	 -53, 	 -50, 	 -50, 	 -61, 	 -79, 	 -46, 	  -4, 	   3, 	  -5, 	 -29, 	 -51, 	   6, 	  23, 	  11, 	  -2, 	 -27, 	 -61, 	 -66, 	 -69, 	 -75, 	 -72, 	 -71, 	 -68, 	 -65, 	 -66, 	 -60, 	 -55, 	 -52, 	 -43, 	 -43, 	
  26, 	  25, 	  29, 	  25, 	  22, 	  21, 	  24, 	  23, 	  21, 	  18, 	  15, 	  18, 	  19, 	  23, 	  24, 	  22, 	  29, 	  25, 	  27, 	  33, 	  33, 	  22, 	  22, 	  15, 	  17, 	  15, 	  24, 	  28, 	  33, 	  46, 	  39, 	  39, 	  42, 	  43, 	  44, 	  48, 	  51, 	  53, 	  53, 	  58, 	  61, 	  64, 	  65, 	  63, 	  68, 	  66, 	  64, 	  64, 	  63, 	  69, 	  65, 	  66, 	  67, 	  63, 	  67, 	  65, 	  65, 	  63, 	  65, 	  64, 	  68, 	  66, 	  67, 	  66, 		  62, 	  61, 	  53, 	  54, 	  58, 	  56, 	  52, 	  50, 	  53, 	  57, 	  53, 	  46, 	  47, 	  45, 	  35, 	  10, 	  -9, 	 -17, 	 -18, 	 -18, 	 -17, 	 -22, 	 -20, 	 -16, 	 -17, 	 -30, 	 -55, 	 -56, 	 -56, 	 -57, 	 -61, 	 -61, 	 -62, 	 -66, 	 -64, 	 -66, 	 -72, 	 -76, 	 -84, 	 -58, 	 -23, 	 -17, 	 -32, 	 -36, 	 -26, 	 -41, 	   6, 	   2, 	   5, 	  -2, 	 -27, 	 -29, 	 -32, 	 -33, 	 -33, 	 -33, 	 -36, 	 -36, 	 -39, 	 -38, 	 -42, 	 -44, 	 -46, 	 -51, 	
  -2, 	  12, 	  10, 	  14, 	  14, 	  18, 	  15, 	  19, 	  18, 	  12, 	   8, 	   8, 	  12, 	  14, 	  18, 	  18, 	  23, 	  20, 	  32, 	  27, 	  29, 	  31, 	  24, 	  28, 	  24, 	  24, 	  21, 	  19, 	  15, 	  17, 	  25, 	  30, 	  36, 	  36, 	  42, 	  45, 	  46, 	  50, 	  48, 	  49, 	  49, 	  50, 	  56, 	  57, 	  62, 	  66, 	  66, 	  67, 	  67, 	  63, 	  64, 	  63, 	  64, 	  66, 	  68, 	  70, 	  68, 	  68, 	  72, 	  72, 	  73, 	  68, 	  70, 	  71, 		  67, 	  63, 	  63, 	  59, 	  59, 	  58, 	  53, 	  47, 	  47, 	  45, 	  46, 	  43, 	  50, 	  49, 	  43, 	  30, 	  15, 	   7, 	 -41, 	 -55, 	 -63, 	 -72, 	 -74, 	 -75, 	 -79, 	 -83, 	 -81, 	 -83, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -84, 	 -84, 	 -87, 	 -87, 	 -85, 	 -83, 	 -59, 	 -33, 	 -36, 	 -35, 	 -34, 	 -25, 	 -53, 	 -37, 	 -35, 	 -48, 	 -42, 	 -60, 	 -63, 	 -66, 	 -66, 	 -67, 	 -66, 	 -72, 	 -63, 	 -69, 	 -67, 	 -69, 	 -74, 	 -64, 	 -76, 	
 -21, 	 -15, 	 -15, 	  -8, 	  -3, 	   1, 	  13, 	  17, 	  22, 	  19, 	  17, 	  17, 	  25, 	  16, 	  17, 	  17, 	  15, 	  15, 	  24, 	  24, 	  26, 	  27, 	  26, 	  24, 	  28, 	  33, 	  31, 	  30, 	  28, 	  20, 	  16, 	   9, 	  13, 	   9, 	  22, 	  30, 	  38, 	  44, 	  54, 	  55, 	  55, 	  49, 	  50, 	  50, 	  47, 	  50, 	  52, 	  60, 	  71, 	  71, 	  70, 	  73, 	  73, 	  76, 	  74, 	  74, 	  75, 	  71, 	  73, 	  72, 	  70, 	  69, 	  66, 	  66, 		  68, 	  64, 	  69, 	  64, 	  65, 	  62, 	  58, 	  55, 	  50, 	  43, 	  36, 	  37, 	  39, 	  41, 	  43, 	  48, 	  35, 	  33, 	   0, 	 -62, 	 -79, 	 -83, 	 -86, 	 -84, 	 -88, 	 -83, 	 -84, 	 -87, 	 -85, 	 -88, 	 -85, 	 -85, 	 -85, 	 -84, 	 -84, 	 -85, 	 -85, 	 -83, 	 -86, 	 -67, 	 -46, 	 -62, 	 -52, 	 -64, 	 -71, 	 -68, 	 -68, 	 -72, 	 -68, 	 -65, 	 -73, 	 -79, 	 -78, 	 -80, 	 -76, 	 -74, 	 -84, 	 -82, 	 -81, 	 -81, 	 -82, 	 -79, 	 -81, 	 -82, 	
 -34, 	 -33, 	 -32, 	 -23, 	 -19, 	 -19, 	 -15, 	  -9, 	  -4, 	   1, 	   8, 	  10, 	  12, 	  10, 	  10, 	  11, 	  13, 	  15, 	  23, 	  25, 	  23, 	  21, 	  20, 	  21, 	  18, 	  25, 	  26, 	  15, 	  21, 	  17, 	  16, 	  16, 	  28, 	  23, 	  10, 	   8, 	  20, 	  35, 	  59, 	  70, 	  78, 	  72, 	  73, 	  58, 	  56, 	  45, 	  47, 	  45, 	  54, 	  80, 	  74, 	  73, 	  72, 	  72, 	  77, 	  72, 	  70, 	  73, 	  69, 	  75, 	  73, 	  67, 	  67, 	  66, 		  67, 	  68, 	  66, 	  70, 	  72, 	  61, 	  62, 	  63, 	  60, 	  54, 	  44, 	  40, 	  42, 	  42, 	  43, 	  48, 	  47, 	  46, 	  33, 	   5, 	 -60, 	 -75, 	 -77, 	 -73, 	 -78, 	 -78, 	 -77, 	 -75, 	 -78, 	 -79, 	 -78, 	 -79, 	 -79, 	 -78, 	 -79, 	 -81, 	 -83, 	 -82, 	 -83, 	 -83, 	 -67, 	 -67, 	 -71, 	 -82, 	 -70, 	 -77, 	 -70, 	 -62, 	 -67, 	 -67, 	 -78, 	 -86, 	 -86, 	 -85, 	 -87, 	 -85, 	 -83, 	 -79, 	 -79, 	 -80, 	 -74, 	 -72, 	 -75, 	 -75, 	
 -45, 	 -46, 	 -40, 	 -40, 	 -35, 	 -30, 	 -29, 	 -27, 	 -22, 	 -18, 	 -16, 	 -10, 	 -10, 	  -4, 	   0, 	   6, 	   4, 	   7, 	   8, 	   8, 	  11, 	  15, 	  17, 	  13, 	  12, 	  10, 	  12, 	   5, 	  10, 	   8, 	  12, 	  14, 	  16, 	  23, 	  20, 	  19, 	  19, 	  26, 	  43, 	  47, 	  58, 	  69, 	  87, 	  87, 	  75, 	  64, 	  55, 	  54, 	  49, 	  45, 	  58, 	  77, 	  81, 	  73, 	  77, 	  70, 	  68, 	  71, 	  67, 	  72, 	  72, 	  76, 	  68, 	  70, 		  68, 	  68, 	  65, 	  63, 	  66, 	  61, 	  63, 	  64, 	  61, 	  63, 	  57, 	  54, 	  47, 	  41, 	  44, 	  48, 	  43, 	  43, 	  46, 	  33, 	   9, 	 -58, 	 -77, 	 -78, 	 -80, 	 -80, 	 -85, 	 -81, 	 -86, 	 -87, 	 -87, 	 -88, 	 -87, 	 -84, 	 -85, 	 -84, 	 -88, 	 -87, 	 -89, 	 -89, 	 -67, 	 -39, 	 -49, 	 -76, 	 -83, 	 -82, 	 -76, 	 -69, 	 -64, 	 -60, 	 -80, 	 -85, 	 -90, 	 -84, 	 -83, 	 -81, 	 -73, 	 -66, 	 -67, 	 -65, 	 -64, 	 -64, 	 -64, 	 -68, 	
 -45, 	 -46, 	 -45, 	 -48, 	 -43, 	 -42, 	 -40, 	 -39, 	 -36, 	 -32, 	 -29, 	 -28, 	 -23, 	 -22, 	 -18, 	 -13, 	 -13, 	  -5, 	  -5, 	  -2, 	  -3, 	  -2, 	   2, 	  -2, 	   0, 	  -1, 	  -2, 	   3, 	   7, 	  13, 	   1, 	   9, 	   4, 	  13, 	  13, 	  19, 	  19, 	  20, 	  15, 	  19, 	  36, 	  53, 	  57, 	  66, 	  86, 	  87, 	  71, 	  49, 	  47, 	  43, 	  65, 	  58, 	  57, 	  79, 	  84, 	  81, 	  72, 	  78, 	  77, 	  71, 	  73, 	  78, 	  67, 	  64, 		  67, 	  67, 	  66, 	  68, 	  63, 	  64, 	  64, 	  63, 	  64, 	  66, 	  64, 	  63, 	  62, 	  55, 	  56, 	  57, 	  55, 	  56, 	  51, 	  42, 	  33, 	   4, 	 -69, 	 -78, 	 -85, 	 -83, 	 -85, 	 -88, 	 -85, 	 -87, 	 -86, 	 -87, 	 -86, 	 -84, 	 -84, 	 -84, 	 -87, 	 -87, 	 -86, 	 -84, 	 -83, 	 -57, 	 -44, 	 -74, 	 -79, 	 -81, 	 -78, 	 -58, 	 -55, 	 -65, 	 -76, 	 -79, 	 -89, 	 -84, 	 -81, 	 -76, 	 -62, 	 -62, 	 -62, 	 -60, 	 -59, 	 -59, 	 -59, 	 -62, 	
 -48, 	 -44, 	 -46, 	 -50, 	 -48, 	 -46, 	 -46, 	 -44, 	 -42, 	 -41, 	 -40, 	 -39, 	 -38, 	 -37, 	 -37, 	 -34, 	 -31, 	 -28, 	 -26, 	 -23, 	 -20, 	 -22, 	 -16, 	 -15, 	 -12, 	 -14, 	 -13, 	  -7, 	  -3, 	  -1, 	  -1, 	  -3, 	  -3, 	   0, 	   1, 	  10, 	   7, 	   5, 	  16, 	   9, 	  12, 	  35, 	  38, 	  30, 	  29, 	  43, 	  55, 	  62, 	  81, 	  76, 	  66, 	  83, 	  55, 	  65, 	  85, 	  85, 	  84, 	  86, 	  83, 	  82, 	  82, 	  75, 	  64, 	  68, 		  61, 	  56, 	  70, 	  62, 	  54, 	  63, 	  61, 	  61, 	  61, 	  61, 	  58, 	  60, 	  63, 	  56, 	  55, 	  56, 	  59, 	  63, 	  62, 	  61, 	  41, 	  43, 	   3, 	 -72, 	 -85, 	 -86, 	 -85, 	 -85, 	 -85, 	 -86, 	 -86, 	 -87, 	 -86, 	 -84, 	 -84, 	 -85, 	 -88, 	 -87, 	 -88, 	 -84, 	 -87, 	 -78, 	 -49, 	 -66, 	 -83, 	 -84, 	 -81, 	 -70, 	 -60, 	 -69, 	 -75, 	 -87, 	 -86, 	 -82, 	 -81, 	 -72, 	 -57, 	 -55, 	 -56, 	 -55, 	 -55, 	 -58, 	 -60, 	 -63, 	
 -48, 	 -46, 	 -47, 	 -46, 	 -44, 	 -44, 	 -47, 	 -41, 	 -47, 	 -47, 	 -44, 	 -47, 	 -46, 	 -49, 	 -48, 	 -44, 	 -45, 	 -45, 	 -40, 	 -42, 	 -37, 	 -37, 	 -36, 	 -30, 	 -24, 	 -25, 	 -21, 	 -15, 	 -14, 	 -11, 	 -12, 	 -10, 	 -12, 	 -11, 	 -11, 	  -2, 	   2, 	  -2, 	   0, 	   5, 	   2, 	   6, 	   2, 	  -7, 	  -2, 	   5, 	  39, 	  51, 	  79, 	  73, 	  69, 	  84, 	  79, 	  32, 	  70, 	  86, 	  88, 	  90, 	  79, 	  87, 	  85, 	  79, 	  73, 	  69, 		  73, 	  55, 	  62, 	  69, 	  60, 	  69, 	  59, 	  64, 	  68, 	  66, 	  61, 	  63, 	  63, 	  63, 	  69, 	  74, 	  69, 	  66, 	  66, 	  65, 	  67, 	  46, 	  43, 	   1, 	 -66, 	 -83, 	 -83, 	 -86, 	 -86, 	 -87, 	 -86, 	 -87, 	 -86, 	 -84, 	 -84, 	 -85, 	 -88, 	 -87, 	 -87, 	 -86, 	 -84, 	 -85, 	 -71, 	 -58, 	 -83, 	 -84, 	 -82, 	 -81, 	 -80, 	 -70, 	 -80, 	 -86, 	 -84, 	 -81, 	 -81, 	 -73, 	 -68, 	 -56, 	 -57, 	 -56, 	 -55, 	 -58, 	 -59, 	 -61, 	
 -51, 	 -49, 	 -53, 	 -48, 	 -46, 	 -47, 	 -43, 	 -43, 	 -42, 	 -46, 	 -48, 	 -49, 	 -52, 	 -55, 	 -54, 	 -56, 	 -55, 	 -54, 	 -53, 	 -53, 	 -54, 	 -54, 	 -47, 	 -45, 	 -42, 	 -39, 	 -38, 	 -31, 	 -27, 	 -22, 	 -17, 	 -14, 	  -8, 	  -6, 	  -8, 	  -5, 	  -4, 	  -6, 	  -5, 	  -7, 	  -3, 	  -3, 	  -7, 	 -15, 	  29, 	   7, 	   9, 	  56, 	  59, 	  81, 	  61, 	  60, 	  78, 	  58, 	  39, 	  59, 	  80, 	  82, 	  93, 	  89, 	  92, 	  71, 	  83, 	  82, 		  88, 	  81, 	  79, 	  81, 	  75, 	  71, 	  73, 	  72, 	  69, 	  68, 	  67, 	  71, 	  73, 	  69, 	  75, 	  71, 	  70, 	  76, 	  73, 	  72, 	  72, 	  65, 	  63, 	  49, 	  20, 	 -67, 	 -81, 	 -83, 	 -85, 	 -85, 	 -86, 	 -88, 	 -86, 	 -86, 	 -86, 	 -87, 	 -88, 	 -89, 	 -87, 	 -87, 	 -87, 	 -89, 	 -83, 	 -79, 	 -83, 	 -82, 	 -76, 	 -77, 	 -72, 	 -67, 	 -78, 	 -85, 	 -82, 	 -79, 	 -80, 	 -71, 	 -67, 	 -65, 	 -59, 	 -59, 	 -56, 	 -61, 	 -63, 	 -63, 	
 -51, 	 -53, 	 -49, 	 -48, 	 -52, 	 -49, 	 -46, 	 -45, 	 -43, 	 -47, 	 -47, 	 -53, 	 -53, 	 -54, 	 -53, 	 -54, 	 -56, 	 -54, 	 -57, 	 -57, 	 -58, 	 -55, 	 -59, 	 -58, 	 -54, 	 -53, 	 -54, 	 -44, 	 -41, 	 -38, 	 -33, 	 -21, 	 -14, 	 -10, 	  -4, 	   0, 	  -4, 	 -10, 	  -9, 	 -10, 	 -13, 	  -9, 	 -11, 	 -11, 	 -14, 	 -23, 	 -21, 	   8, 	  47, 	  36, 	  68, 	  89, 	  88, 	  82, 	  38, 	  23, 	  57, 	  82, 	  88, 	  95, 	  92, 	  87, 	  82, 	  84, 		  90, 	  86, 	  88, 	  85, 	  83, 	  80, 	  75, 	  71, 	  76, 	  72, 	  70, 	  67, 	  70, 	  67, 	  72, 	  71, 	  74, 	  70, 	  76, 	  73, 	  77, 	  78, 	  75, 	  59, 	  49, 	   6, 	 -78, 	 -83, 	 -85, 	 -86, 	 -87, 	 -88, 	 -88, 	 -87, 	 -87, 	 -88, 	 -88, 	 -90, 	 -91, 	 -87, 	 -86, 	 -84, 	 -85, 	 -82, 	 -84, 	 -80, 	 -80, 	 -79, 	 -75, 	 -65, 	 -75, 	 -84, 	 -82, 	 -82, 	 -81, 	 -69, 	 -71, 	 -63, 	 -61, 	 -61, 	 -62, 	 -62, 	 -59, 	 -59, 	
 -50, 	 -53, 	 -50, 	 -46, 	 -46, 	 -52, 	 -49, 	 -49, 	 -48, 	 -47, 	 -50, 	 -53, 	 -53, 	 -53, 	 -54, 	 -55, 	 -53, 	 -54, 	 -55, 	 -58, 	 -59, 	 -61, 	 -62, 	 -62, 	 -52, 	 -57, 	 -64, 	 -58, 	 -55, 	 -52, 	 -38, 	 -30, 	 -25, 	 -16, 	 -14, 	  -8, 	  -6, 	  -9, 	  -8, 	  -4, 	  -8, 	 -12, 	 -12, 	 -10, 	 -15, 	 -21, 	 -25, 	 -17, 	  43, 	  27, 	   9, 	  53, 	  80, 	  89, 	  80, 	  38, 	  16, 	  42, 	  75, 	  89, 	  92, 	  88, 	  90, 	  92, 		  92, 	  92, 	  89, 	  89, 	  86, 	  86, 	  80, 	  78, 	  75, 	  75, 	  75, 	  71, 	  73, 	  74, 	  76, 	  77, 	  78, 	  79, 	  78, 	  72, 	  72, 	  78, 	  79, 	  74, 	  59, 	  44, 	 -14, 	 -80, 	 -83, 	 -86, 	 -86, 	 -88, 	 -87, 	 -86, 	 -86, 	 -86, 	 -87, 	 -88, 	 -88, 	 -83, 	 -86, 	 -82, 	 -83, 	 -84, 	 -80, 	 -80, 	 -80, 	 -77, 	 -74, 	 -66, 	 -72, 	 -81, 	 -82, 	 -83, 	 -78, 	 -71, 	 -70, 	 -67, 	 -58, 	 -59, 	 -60, 	 -60, 	 -58, 	 -63, 	
 -45, 	 -42, 	 -39, 	 -39, 	 -40, 	 -44, 	 -46, 	 -49, 	 -47, 	 -46, 	 -49, 	 -52, 	 -50, 	 -54, 	 -56, 	 -54, 	 -57, 	 -53, 	 -54, 	 -58, 	 -59, 	 -58, 	 -62, 	 -62, 	 -62, 	 -63, 	 -64, 	 -66, 	 -65, 	 -61, 	 -51, 	 -43, 	 -33, 	 -26, 	 -17, 	 -13, 	  -9, 	  -5, 	 -10, 	  -7, 	  -7, 	  -9, 	 -10, 	  -5, 	 -10, 	 -17, 	 -23, 	 -29, 	 -28, 	   0, 	  29, 	   2, 	  28, 	  71, 	  79, 	  72, 	  25, 	   1, 	  13, 	  71, 	  90, 	  92, 	  92, 	  94, 		  95, 	  95, 	  89, 	  88, 	  85, 	  88, 	  83, 	  81, 	  81, 	  83, 	  76, 	  79, 	  76, 	  75, 	  77, 	  80, 	  81, 	  79, 	  83, 	  78, 	  71, 	  74, 	  76, 	  76, 	  71, 	  57, 	  47, 	 -26, 	 -78, 	 -85, 	 -85, 	 -87, 	 -86, 	 -84, 	 -84, 	 -85, 	 -84, 	 -89, 	 -85, 	 -85, 	 -85, 	 -81, 	 -83, 	 -83, 	 -81, 	 -80, 	 -80, 	 -74, 	 -73, 	 -66, 	 -69, 	 -82, 	 -80, 	 -82, 	 -76, 	 -73, 	 -68, 	 -65, 	 -61, 	 -61, 	 -59, 	 -57, 	 -59, 	 -55, 	
 -72, 	 -71, 	 -66, 	 -59, 	 -52, 	 -45, 	 -42, 	 -37, 	 -34, 	 -39, 	 -48, 	 -50, 	 -53, 	 -56, 	 -59, 	 -59, 	 -59, 	 -58, 	 -59, 	 -59, 	 -60, 	 -64, 	 -63, 	 -63, 	 -62, 	 -63, 	 -67, 	 -63, 	 -67, 	 -68, 	 -62, 	 -56, 	 -45, 	 -34, 	 -24, 	 -15, 	 -13, 	  -7, 	 -11, 	 -10, 	  -7, 	  -6, 	  -3, 	  -6, 	  -8, 	 -15, 	 -20, 	 -25, 	 -34, 	 -33, 	 -20, 	 -19, 	 -11, 	   7, 	  18, 	  54, 	  59, 	  26, 	   3, 	  22, 	  76, 	  87, 	  92, 	  88, 		  92, 	  94, 	  90, 	  92, 	  90, 	  91, 	  90, 	  85, 	  86, 	  84, 	  81, 	  83, 	  79, 	  80, 	  79, 	  80, 	  83, 	  83, 	  79, 	  81, 	  81, 	  81, 	  81, 	  78, 	  76, 	  67, 	  51, 	  51, 	 -43, 	 -80, 	 -79, 	 -82, 	 -80, 	 -84, 	 -78, 	 -83, 	 -84, 	 -85, 	 -85, 	 -84, 	 -82, 	 -81, 	 -82, 	 -82, 	 -82, 	 -79, 	 -77, 	 -74, 	 -78, 	 -69, 	 -67, 	 -81, 	 -83, 	 -82, 	 -75, 	 -70, 	 -68, 	 -61, 	 -61, 	 -58, 	 -56, 	 -57, 	 -55, 	 -49, 	
 -79, 	 -78, 	 -75, 	 -75, 	 -75, 	 -72, 	 -72, 	 -69, 	 -61, 	 -54, 	 -48, 	 -41, 	 -48, 	 -52, 	 -58, 	 -59, 	 -66, 	 -62, 	 -60, 	 -59, 	 -60, 	 -62, 	 -62, 	 -63, 	 -66, 	 -67, 	 -64, 	 -65, 	 -68, 	 -68, 	 -68, 	 -64, 	 -59, 	 -47, 	 -32, 	 -24, 	 -17, 	 -11, 	 -13, 	 -15, 	 -11, 	  -6, 	  -5, 	 -10, 	  -6, 	 -14, 	 -15, 	 -22, 	 -28, 	 -39, 	 -36, 	 -33, 	 -28, 	 -18, 	 -16, 	  -6, 	  21, 	  66, 	  20, 	  -3, 	  24, 	  77, 	  89, 	  90, 		  92, 	  91, 	  90, 	  92, 	  92, 	  92, 	  89, 	  88, 	  83, 	  86, 	  82, 	  78, 	  65, 	  78, 	  81, 	  82, 	  81, 	  81, 	  84, 	  81, 	  77, 	  81, 	  83, 	  84, 	  79, 	  78, 	  61, 	  60, 	  37, 	 -68, 	 -75, 	 -80, 	 -79, 	 -83, 	 -82, 	 -81, 	 -84, 	 -84, 	 -85, 	 -83, 	 -81, 	 -81, 	 -80, 	 -79, 	 -81, 	 -79, 	 -77, 	 -79, 	 -78, 	 -68, 	 -67, 	 -83, 	 -86, 	 -82, 	 -62, 	 -51, 	 -40, 	 -42, 	 -49, 	 -53, 	 -53, 	 -43, 	 -30, 	 -17, 	
 -81, 	 -79, 	 -81, 	 -79, 	 -80, 	 -79, 	 -80, 	 -79, 	 -78, 	 -75, 	 -76, 	 -70, 	 -57, 	 -49, 	 -50, 	 -55, 	 -60, 	 -59, 	 -59, 	 -64, 	 -66, 	 -63, 	 -62, 	 -61, 	 -61, 	 -61, 	 -67, 	 -62, 	 -67, 	 -68, 	 -67, 	 -66, 	 -68, 	 -58, 	 -47, 	 -33, 	 -18, 	 -10, 	 -15, 	 -13, 	 -17, 	 -12, 	  -7, 	 -13, 	  -7, 	 -13, 	 -13, 	 -15, 	 -27, 	 -32, 	 -39, 	 -38, 	 -35, 	 -28, 	 -28, 	 -21, 	 -12, 	  43, 	  49, 	 -17, 	  -9, 	  33, 	  81, 	  91, 		  89, 	  92, 	  74, 	  83, 	  72, 	  72, 	  79, 	  83, 	  76, 	  66, 	  77, 	  77, 	  69, 	  72, 	  74, 	  83, 	  78, 	  63, 	  80, 	  82, 	  82, 	  82, 	  86, 	  83, 	  84, 	  81, 	  76, 	  59, 	  67, 	  -1, 	 -75, 	 -74, 	 -79, 	 -80, 	 -81, 	 -78, 	 -84, 	 -83, 	 -86, 	 -85, 	 -83, 	 -83, 	 -82, 	 -81, 	 -80, 	 -81, 	 -81, 	 -81, 	 -78, 	 -68, 	 -68, 	 -85, 	 -86, 	 -81, 	 -63, 	 -47, 	 -22, 	 -17, 	 -12, 	 -20, 	 -28, 	 -22, 	 -12, 	  17, 	
 -80, 	 -79, 	 -79, 	 -80, 	 -79, 	 -77, 	 -79, 	 -80, 	 -77, 	 -77, 	 -78, 	 -76, 	 -76, 	 -73, 	 -63, 	 -49, 	 -42, 	 -51, 	 -60, 	 -59, 	 -62, 	 -65, 	 -62, 	 -62, 	 -62, 	 -62, 	 -63, 	 -68, 	 -64, 	 -65, 	 -67, 	 -66, 	 -67, 	 -65, 	 -57, 	 -45, 	 -25, 	 -17, 	 -18, 	 -26, 	 -23, 	 -20, 	 -14, 	 -13, 	 -13, 	  -8, 	 -13, 	 -19, 	 -21, 	 -25, 	 -39, 	 -40, 	 -42, 	 -30, 	 -37, 	 -29, 	 -25, 	 -17, 	  -1, 	   7, 	 -24, 	  -9, 	  52, 	  82, 		  87, 	  84, 	  75, 	  65, 	  61, 	  64, 	  74, 	  81, 	  76, 	  67, 	  71, 	  69, 	  71, 	  75, 	  77, 	  76, 	  65, 	  50, 	  64, 	  85, 	  81, 	  76, 	  73, 	  86, 	  84, 	  83, 	  78, 	  72, 	  68, 	  54, 	 -50, 	 -75, 	 -76, 	 -78, 	 -79, 	 -80, 	 -82, 	 -82, 	 -83, 	 -82, 	 -80, 	 -83, 	 -83, 	 -80, 	 -80, 	 -82, 	 -84, 	 -82, 	 -78, 	 -71, 	 -68, 	 -84, 	 -89, 	 -77, 	 -62, 	 -46, 	 -32, 	 -24, 	 -22, 	 -21, 	 -22, 	 -16, 	   0, 	  63, 	
 -85, 	 -83, 	 -81, 	 -81, 	 -80, 	 -79, 	 -82, 	 -79, 	 -81, 	 -80, 	 -81, 	 -79, 	 -79, 	 -76, 	 -76, 	 -74, 	 -61, 	 -46, 	 -44, 	 -55, 	 -60, 	 -60, 	 -63, 	 -59, 	 -64, 	 -61, 	 -63, 	 -65, 	 -63, 	 -64, 	 -63, 	 -64, 	 -68, 	 -68, 	 -67, 	 -56, 	 -45, 	 -28, 	 -21, 	 -28, 	 -26, 	 -24, 	 -20, 	 -15, 	 -13, 	 -18, 	 -17, 	 -19, 	 -22, 	 -21, 	 -29, 	 -45, 	 -46, 	 -39, 	 -41, 	 -41, 	 -36, 	 -34, 	 -24, 	 -21, 	 -27, 	 -23, 	   3, 	  58, 		  64, 	  65, 	  78, 	  78, 	  75, 	  73, 	  72, 	  74, 	  69, 	  73, 	  74, 	  72, 	  73, 	  66, 	  70, 	  71, 	  70, 	  59, 	  58, 	  67, 	  68, 	  71, 	  56, 	  78, 	  75, 	  76, 	  72, 	  79, 	  65, 	  61, 	  19, 	 -72, 	 -75, 	 -76, 	 -79, 	 -81, 	 -81, 	 -83, 	 -81, 	 -80, 	 -84, 	 -83, 	 -79, 	 -80, 	 -79, 	 -82, 	 -84, 	 -80, 	 -80, 	 -73, 	 -64, 	 -86, 	 -85, 	 -75, 	 -62, 	 -56, 	 -53, 	 -38, 	 -32, 	 -25, 	 -27, 	  -9, 	  51, 	  68, 	
 -93, 	 -94, 	 -91, 	 -90, 	 -89, 	 -85, 	 -84, 	 -82, 	 -81, 	 -81, 	 -81, 	 -82, 	 -80, 	 -79, 	 -78, 	 -76, 	 -77, 	 -70, 	 -52, 	 -38, 	 -49, 	 -59, 	 -63, 	 -58, 	 -59, 	 -62, 	 -59, 	 -63, 	 -65, 	 -62, 	 -62, 	 -63, 	 -68, 	 -68, 	 -68, 	 -64, 	 -56, 	 -42, 	 -22, 	 -13, 	 -20, 	 -17, 	 -18, 	 -20, 	 -20, 	 -16, 	 -19, 	 -20, 	 -17, 	 -20, 	 -27, 	 -37, 	 -50, 	 -47, 	 -53, 	 -44, 	 -45, 	 -39, 	 -36, 	 -31, 	 -33, 	 -25, 	 -17, 	  40, 		  72, 	  75, 	  79, 	  71, 	  68, 	  78, 	  72, 	  68, 	  66, 	  66, 	  66, 	  66, 	  73, 	  64, 	  61, 	  67, 	  69, 	  67, 	  63, 	  49, 	  44, 	  58, 	  50, 	  55, 	  69, 	  73, 	  58, 	  80, 	  72, 	  64, 	  52, 	 -35, 	 -72, 	 -76, 	 -79, 	 -79, 	 -78, 	 -80, 	 -81, 	 -82, 	 -81, 	 -80, 	 -79, 	 -80, 	 -81, 	 -81, 	 -81, 	 -79, 	 -81, 	 -74, 	 -63, 	 -82, 	 -84, 	 -75, 	 -64, 	 -58, 	 -66, 	 -52, 	 -38, 	 -35, 	 -21, 	  23, 	  74, 	  13, 	
 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -91, 	 -91, 	 -87, 	 -85, 	 -83, 	 -80, 	 -79, 	 -79, 	 -78, 	 -78, 	 -75, 	 -70, 	 -59, 	 -40, 	 -44, 	 -56, 	 -60, 	 -63, 	 -59, 	 -61, 	 -66, 	 -67, 	 -65, 	 -65, 	 -66, 	 -67, 	 -67, 	 -68, 	 -66, 	 -63, 	 -50, 	 -31, 	  -5, 	 -14, 	 -21, 	 -21, 	 -17, 	 -25, 	 -22, 	 -26, 	 -29, 	 -23, 	 -20, 	 -26, 	 -30, 	 -47, 	 -44, 	 -48, 	 -51, 	 -47, 	 -42, 	 -42, 	 -43, 	 -33, 	 -32, 	  36, 	  61, 		  67, 	  68, 	  70, 	  66, 	  64, 	  64, 	  65, 	  72, 	  68, 	  60, 	  65, 	  66, 	  61, 	  61, 	  61, 	  59, 	  64, 	  61, 	  63, 	  62, 	  59, 	  56, 	  49, 	  45, 	  51, 	  61, 	  58, 	  62, 	  79, 	  68, 	  59, 	  18, 	 -62, 	 -66, 	 -67, 	 -64, 	 -69, 	 -72, 	 -78, 	 -84, 	 -78, 	 -75, 	 -80, 	 -83, 	 -83, 	 -80, 	 -78, 	 -81, 	 -81, 	 -77, 	 -60, 	 -82, 	 -79, 	 -65, 	 -53, 	 -41, 	 -63, 	 -68, 	 -54, 	 -48, 	 -17, 	  56, 	  46, 	 -35, 	
 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -96, 	 -93, 	 -90, 	 -93, 	 -92, 	 -88, 	 -85, 	 -80, 	 -78, 	 -81, 	 -78, 	 -74, 	 -76, 	 -62, 	 -40, 	 -41, 	 -56, 	 -63, 	 -60, 	 -61, 	 -65, 	 -66, 	 -68, 	 -65, 	 -66, 	 -68, 	 -68, 	 -66, 	 -66, 	 -68, 	 -61, 	 -48, 	 -16, 	  14, 	 -19, 	 -27, 	 -28, 	 -33, 	 -32, 	 -26, 	 -34, 	 -30, 	 -30, 	 -26, 	 -26, 	 -40, 	 -51, 	 -52, 	 -50, 	 -51, 	 -45, 	 -47, 	 -49, 	 -40, 	  -9, 	  72, 	  78, 		  78, 	  76, 	  77, 	  75, 	  75, 	  73, 	  69, 	  71, 	  68, 	  65, 	  70, 	  73, 	  67, 	  66, 	  68, 	  66, 	  64, 	  63, 	  64, 	  62, 	  67, 	  62, 	  56, 	  51, 	  47, 	  47, 	  58, 	  51, 	  75, 	  75, 	  59, 	  50, 	 -29, 	 -46, 	 -53, 	 -56, 	 -56, 	 -66, 	 -69, 	 -75, 	 -80, 	 -80, 	 -80, 	 -83, 	 -82, 	 -77, 	 -72, 	 -69, 	 -79, 	 -77, 	 -60, 	 -79, 	 -78, 	 -67, 	 -63, 	 -47, 	 -46, 	 -57, 	 -60, 	 -40, 	  41, 	  63, 	  -5, 	 -14, 	
 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -93, 	 -93, 	 -93, 	 -93, 	 -92, 	 -91, 	 -88, 	 -83, 	 -79, 	 -79, 	 -79, 	 -77, 	 -76, 	 -72, 	 -45, 	 -36, 	 -60, 	 -61, 	 -61, 	 -64, 	 -64, 	 -68, 	 -67, 	 -67, 	 -68, 	 -68, 	 -66, 	 -66, 	 -68, 	 -69, 	 -54, 	 -32, 	  36, 	  13, 	 -30, 	 -30, 	 -28, 	 -35, 	 -34, 	 -37, 	 -34, 	 -34, 	 -33, 	 -29, 	 -35, 	 -27, 	 -53, 	 -53, 	 -53, 	 -49, 	 -51, 	 -52, 	 -41, 	  20, 	  60, 	  73, 		  72, 	  77, 	  78, 	  73, 	  74, 	  72, 	  75, 	  76, 	  74, 	  76, 	  77, 	  74, 	  79, 	  80, 	  80, 	  78, 	  75, 	  78, 	  79, 	  79, 	  77, 	  81, 	  78, 	  76, 	  75, 	  71, 	  67, 	  61, 	  70, 	  67, 	  51, 	  46, 	  12, 	 -53, 	 -57, 	 -54, 	 -54, 	 -53, 	 -59, 	 -67, 	 -79, 	 -84, 	 -84, 	 -83, 	 -82, 	 -79, 	 -72, 	 -68, 	 -78, 	 -78, 	 -61, 	 -77, 	 -77, 	 -68, 	 -68, 	 -61, 	 -59, 	 -66, 	 -52, 	  13, 	  70, 	  25, 	 -16, 	 -13, 	
 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -93, 	 -93, 	 -93, 	 -94, 	 -92, 	 -92, 	 -91, 	 -88, 	 -81, 	 -77, 	 -76, 	 -78, 	 -76, 	 -71, 	 -44, 	 -37, 	 -54, 	 -63, 	 -66, 	 -66, 	 -64, 	 -68, 	 -68, 	 -68, 	 -68, 	 -65, 	 -66, 	 -67, 	 -68, 	 -59, 	 -45, 	   2, 	  66, 	  -5, 	 -28, 	 -28, 	 -33, 	 -42, 	 -39, 	 -36, 	 -35, 	 -31, 	 -28, 	 -29, 	 -41, 	 -57, 	 -55, 	 -55, 	 -56, 	 -54, 	 -52, 	 -28, 	  28, 	  25, 	   4, 		  -1, 	   7, 	   9, 	  14, 	  20, 	  25, 	  33, 	  39, 	  46, 	  53, 	  55, 	  57, 	  61, 	  60, 	  55, 	  58, 	  64, 	  66, 	  66, 	  64, 	  64, 	  64, 	  55, 	  45, 	  34, 	  20, 	   3, 	  -6, 	 -14, 	 -21, 	 -38, 	 -48, 	 -50, 	 -62, 	 -61, 	 -61, 	 -63, 	 -58, 	 -60, 	 -67, 	 -79, 	 -83, 	 -85, 	 -83, 	 -83, 	 -79, 	 -76, 	 -73, 	 -86, 	 -75, 	 -62, 	 -73, 	 -68, 	 -59, 	 -56, 	 -54, 	 -47, 	 -52, 	 -12, 	  62, 	  47, 	 -11, 	 -15, 	 -19, 	
 -92, 	 -92, 	 -93, 	 -93, 	 -93, 	 -93, 	 -94, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -87, 	 -83, 	 -78, 	 -79, 	 -79, 	 -77, 	 -70, 	 -44, 	 -35, 	 -59, 	 -64, 	 -64, 	 -69, 	 -67, 	 -66, 	 -67, 	 -67, 	 -62, 	 -69, 	 -68, 	 -66, 	 -66, 	 -52, 	 -27, 	  64, 	  39, 	 -19, 	 -28, 	 -28, 	 -34, 	 -38, 	 -37, 	 -39, 	 -38, 	 -34, 	 -31, 	 -40, 	 -55, 	 -59, 	 -58, 	 -59, 	 -61, 	 -56, 	 -36, 	   3, 	 -27, 	 -29, 		 -15, 	 -25, 	 -49, 	 -58, 	 -60, 	 -51, 	 -41, 	 -27, 	 -18, 	 -12, 	 -19, 	 -31, 	 -39, 	 -36, 	 -32, 	 -34, 	 -31, 	 -43, 	 -53, 	 -51, 	 -53, 	 -58, 	 -56, 	 -50, 	 -56, 	 -65, 	 -69, 	 -76, 	 -74, 	 -78, 	 -76, 	 -82, 	 -83, 	 -77, 	 -68, 	 -66, 	 -70, 	 -68, 	 -69, 	 -76, 	 -80, 	 -83, 	 -85, 	 -83, 	 -85, 	 -81, 	 -77, 	 -78, 	 -80, 	 -75, 	 -58, 	 -68, 	 -47, 	 -38, 	 -37, 	 -25, 	 -20, 	  -3, 	  55, 	  58, 	 -10, 	 -31, 	 -30, 	 -24, 	
 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -92, 	 -91, 	 -91, 	 -86, 	 -81, 	 -78, 	 -81, 	 -73, 	 -70, 	 -44, 	 -38, 	 -57, 	 -59, 	 -65, 	 -65, 	 -66, 	 -66, 	 -68, 	 -65, 	 -67, 	 -66, 	 -66, 	 -62, 	 -58, 	 -45, 	  41, 	  80, 	  -9, 	 -29, 	 -28, 	 -30, 	 -38, 	 -39, 	 -42, 	 -44, 	 -40, 	 -39, 	 -42, 	 -53, 	 -60, 	 -63, 	 -61, 	 -62, 	 -61, 	 -57, 	 -28, 	 -77, 	 -74, 		 -66, 	 -52, 	 -61, 	 -68, 	 -66, 	 -50, 	 -48, 	 -44, 	 -65, 	 -61, 	 -52, 	 -75, 	 -74, 	 -73, 	 -66, 	 -71, 	 -57, 	 -54, 	 -42, 	 -39, 	 -36, 	 -40, 	 -28, 	 -20, 	 -20, 	 -22, 	 -28, 	 -45, 	 -75, 	 -77, 	 -84, 	 -86, 	 -86, 	 -79, 	 -67, 	 -73, 	 -73, 	 -71, 	 -79, 	 -83, 	 -84, 	 -83, 	 -84, 	 -84, 	 -84, 	 -81, 	 -78, 	 -83, 	 -82, 	 -74, 	 -57, 	 -66, 	 -48, 	 -36, 	 -44, 	 -49, 	 -41, 	  13, 	  70, 	   3, 	 -44, 	 -47, 	 -22, 	 -23, 	
 -91, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -93, 	 -94, 	 -93, 	 -92, 	 -91, 	 -85, 	 -79, 	 -80, 	 -78, 	 -76, 	 -69, 	 -31, 	 -41, 	 -56, 	 -61, 	 -63, 	 -65, 	 -68, 	 -68, 	 -68, 	 -65, 	 -69, 	 -69, 	 -66, 	 -64, 	 -51, 	   0, 	  80, 	  17, 	 -18, 	 -31, 	 -37, 	 -37, 	 -37, 	 -39, 	 -38, 	 -39, 	 -37, 	 -39, 	 -48, 	 -60, 	 -60, 	 -64, 	 -61, 	 -65, 	 -64, 	 -33, 	 -63, 	 -69, 		 -50, 	 -64, 	 -62, 	 -70, 	 -73, 	 -59, 	 -40, 	 -37, 	 -68, 	 -71, 	 -69, 	 -55, 	 -49, 	 -66, 	 -80, 	 -27, 	  -8, 	 -11, 	 -25, 	 -37, 	 -48, 	 -55, 	 -54, 	 -53, 	 -50, 	 -43, 	 -46, 	 -58, 	 -65, 	 -77, 	 -81, 	 -82, 	 -83, 	 -74, 	 -61, 	 -66, 	 -67, 	 -71, 	 -79, 	 -84, 	 -82, 	 -81, 	 -84, 	 -85, 	 -83, 	 -79, 	 -68, 	 -79, 	 -82, 	 -74, 	 -50, 	 -54, 	 -55, 	 -51, 	 -54, 	 -51, 	 -19, 	  59, 	  39, 	 -12, 	 -20, 	 -18, 	 -16, 	 -23, 	
 -92, 	 -90, 	 -90, 	 -93, 	 -91, 	 -91, 	 -93, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -92, 	 -92, 	 -87, 	 -80, 	 -78, 	 -78, 	 -76, 	 -61, 	 -29, 	 -47, 	 -60, 	 -60, 	 -63, 	 -67, 	 -68, 	 -65, 	 -65, 	 -66, 	 -69, 	 -67, 	 -65, 	 -55, 	 -25, 	  54, 	  47, 	 -11, 	 -29, 	 -35, 	 -41, 	 -38, 	 -36, 	 -34, 	 -36, 	 -38, 	 -30, 	 -46, 	 -58, 	 -62, 	 -59, 	 -62, 	 -65, 	 -67, 	 -43, 	  -5, 	 -39, 		 -37, 	 -42, 	 -71, 	 -71, 	 -74, 	 -68, 	 -52, 	 -50, 	 -65, 	 -71, 	 -59, 	  -4, 	  36, 	  -9, 	 -70, 	 -47, 	 -38, 	 -49, 	 -63, 	 -66, 	 -69, 	 -73, 	 -73, 	 -68, 	 -59, 	 -50, 	 -52, 	 -64, 	 -63, 	 -66, 	 -61, 	 -44, 	 -74, 	 -63, 	   9, 	 -35, 	 -69, 	 -74, 	 -73, 	 -76, 	 -82, 	 -83, 	 -84, 	 -86, 	 -81, 	 -77, 	 -70, 	 -76, 	 -79, 	 -74, 	 -53, 	 -42, 	 -46, 	 -54, 	 -52, 	 -38, 	   3, 	  33, 	 -22, 	 -24, 	 -22, 	 -24, 	 -30, 	 -44, 	
 -89, 	 -89, 	 -91, 	 -93, 	 -92, 	 -90, 	 -93, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -90, 	 -86, 	 -81, 	 -76, 	 -77, 	 -74, 	 -57, 	 -29, 	 -50, 	 -58, 	 -62, 	 -64, 	 -67, 	 -68, 	 -64, 	 -69, 	 -71, 	 -70, 	 -64, 	 -60, 	 -42, 	  16, 	  76, 	   8, 	 -26, 	 -35, 	 -41, 	 -42, 	 -39, 	 -35, 	 -35, 	 -34, 	 -36, 	 -39, 	 -51, 	 -64, 	 -63, 	 -64, 	 -68, 	 -70, 	 -63, 	   2, 	 -35, 		 -28, 	 -58, 	 -73, 	 -72, 	 -75, 	 -69, 	 -52, 	 -56, 	 -60, 	 -71, 	 -60, 	 -22, 	  45, 	  17, 	 -59, 	 -51, 	 -37, 	 -50, 	 -60, 	 -62, 	 -66, 	 -69, 	 -73, 	 -72, 	 -73, 	 -50, 	 -49, 	 -62, 	 -71, 	 -32, 	   7, 	   2, 	 -73, 	 -57, 	  12, 	 -18, 	 -65, 	 -78, 	 -78, 	 -73, 	 -73, 	 -75, 	 -80, 	 -80, 	 -79, 	 -76, 	 -72, 	 -85, 	 -82, 	 -77, 	 -54, 	 -43, 	 -49, 	 -45, 	 -36, 	 -18, 	  -9, 	 -35, 	 -49, 	 -48, 	 -40, 	 -38, 	 -55, 	 -68, 	
 -89, 	 -88, 	 -90, 	 -92, 	 -92, 	 -90, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -90, 	 -91, 	 -92, 	 -92, 	 -92, 	 -93, 	 -86, 	 -80, 	 -78, 	 -75, 	 -75, 	 -49, 	 -30, 	 -53, 	 -60, 	 -64, 	 -71, 	 -68, 	 -70, 	 -70, 	 -67, 	 -72, 	 -66, 	 -63, 	 -52, 	 -14, 	  66, 	  39, 	 -18, 	 -29, 	 -37, 	 -40, 	 -34, 	 -32, 	 -37, 	 -32, 	 -34, 	 -41, 	 -40, 	 -58, 	 -63, 	 -64, 	 -64, 	 -66, 	 -72, 	 -28, 	 -45, 		 -72, 	 -76, 	 -77, 	 -72, 	 -72, 	 -68, 	 -61, 	 -48, 	 -61, 	 -69, 	 -68, 	 -51, 	  16, 	  -2, 	 -62, 	 -52, 	 -46, 	 -52, 	 -59, 	 -58, 	 -66, 	 -70, 	 -74, 	 -77, 	 -77, 	 -73, 	 -67, 	 -70, 	 -65, 	 -51, 	 -17, 	 -54, 	 -72, 	 -58, 	  26, 	 -37, 	 -68, 	 -78, 	 -79, 	 -80, 	 -75, 	 -73, 	 -65, 	 -61, 	 -67, 	 -70, 	 -72, 	 -72, 	 -81, 	 -76, 	 -59, 	 -52, 	 -51, 	 -35, 	   2, 	  61, 	 -13, 	 -44, 	 -47, 	 -44, 	 -51, 	 -58, 	 -63, 	 -67, 	
 -89, 	 -89, 	 -90, 	 -89, 	 -90, 	 -89, 	 -90, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -87, 	 -78, 	 -77, 	 -77, 	 -71, 	 -40, 	 -38, 	 -55, 	 -60, 	 -69, 	 -68, 	 -68, 	 -71, 	 -69, 	 -71, 	 -67, 	 -65, 	 -61, 	 -37, 	  34, 	  73, 	  -5, 	 -30, 	 -39, 	 -34, 	 -29, 	 -30, 	 -36, 	 -36, 	 -33, 	 -36, 	 -34, 	 -47, 	 -62, 	 -61, 	 -63, 	 -60, 	 -68, 	 -61, 	 -21, 		 -70, 	 -82, 	 -79, 	 -66, 	 -55, 	 -62, 	 -70, 	 -70, 	 -62, 	 -69, 	 -73, 	 -71, 	 -58, 	 -62, 	 -63, 	 -55, 	 -50, 	 -52, 	 -51, 	 -55, 	 -58, 	 -68, 	 -66, 	 -67, 	 -65, 	 -77, 	 -78, 	 -71, 	 -52, 	  10, 	 -36, 	 -69, 	 -74, 	 -59, 	  35, 	   2, 	 -70, 	 -76, 	 -77, 	 -80, 	 -81, 	 -77, 	 -58, 	 -62, 	 -74, 	 -69, 	 -74, 	 -77, 	 -81, 	 -77, 	 -59, 	 -45, 	 -49, 	 -21, 	  59, 	  57, 	 -28, 	 -46, 	 -34, 	 -36, 	 -49, 	 -63, 	 -66, 	 -72, 	
 -82, 	 -88, 	 -87, 	 -91, 	 -90, 	 -90, 	 -88, 	 -91, 	 -91, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -92, 	 -92, 	 -91, 	 -92, 	 -94, 	 -93, 	 -89, 	 -83, 	 -80, 	 -78, 	 -75, 	 -69, 	 -33, 	 -46, 	 -58, 	 -66, 	 -66, 	 -69, 	 -67, 	 -67, 	 -67, 	 -66, 	 -62, 	 -61, 	 -49, 	  -2, 	  78, 	  19, 	 -23, 	 -35, 	 -33, 	 -28, 	 -33, 	 -30, 	 -36, 	 -39, 	 -38, 	 -38, 	 -40, 	 -62, 	 -61, 	 -63, 	 -63, 	 -64, 	 -63, 	 -25, 		 -66, 	 -70, 	 -74, 	 -76, 	 -67, 	 -63, 	 -62, 	 -71, 	 -65, 	 -55, 	 -57, 	 -41, 	 -60, 	 -73, 	 -59, 	 -54, 	 -50, 	 -52, 	 -55, 	 -61, 	 -45, 	 -69, 	 -66, 	 -68, 	 -63, 	 -78, 	 -78, 	 -78, 	 -45, 	 -52, 	 -75, 	 -75, 	 -77, 	 -54, 	  33, 	  35, 	 -57, 	 -68, 	 -74, 	 -79, 	 -80, 	 -76, 	 -45, 	 -39, 	 -69, 	 -70, 	 -75, 	 -78, 	 -81, 	 -70, 	 -56, 	 -34, 	 -25, 	  34, 	  71, 	   2, 	 -39, 	 -42, 	 -38, 	 -50, 	 -59, 	 -65, 	 -66, 	 -74, 	
 -80, 	 -87, 	 -87, 	 -89, 	 -87, 	 -87, 	 -87, 	 -89, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -91, 	 -90, 	 -91, 	 -93, 	 -93, 	 -93, 	 -89, 	 -83, 	 -78, 	 -79, 	 -75, 	 -62, 	 -32, 	 -50, 	 -61, 	 -64, 	 -67, 	 -70, 	 -72, 	 -70, 	 -67, 	 -65, 	 -65, 	 -56, 	 -29, 	  45, 	  51, 	 -18, 	 -32, 	 -29, 	 -35, 	 -33, 	 -31, 	 -31, 	 -32, 	 -34, 	 -38, 	 -38, 	 -52, 	 -64, 	 -61, 	 -65, 	 -68, 	 -69, 	 -43, 		 -10, 	 -25, 	 -70, 	 -74, 	 -72, 	 -67, 	 -67, 	 -73, 	 -66, 	 -53, 	 -37, 	  -6, 	   5, 	 -43, 	 -74, 	 -66, 	 -61, 	 -65, 	 -70, 	 -72, 	 -76, 	 -80, 	 -76, 	 -80, 	 -84, 	 -83, 	 -86, 	 -84, 	 -74, 	 -66, 	 -73, 	 -65, 	 -74, 	 -48, 	  43, 	  45, 	 -29, 	 -70, 	 -77, 	 -75, 	 -82, 	 -83, 	 -75, 	 -70, 	 -71, 	 -71, 	 -73, 	 -79, 	 -76, 	 -78, 	 -62, 	 -38, 	  -7, 	  65, 	  34, 	 -28, 	 -38, 	 -36, 	 -47, 	 -57, 	 -63, 	 -65, 	 -69, 	 -75, 	
 -75, 	 -81, 	 -84, 	 -86, 	 -86, 	 -86, 	 -88, 	 -87, 	 -86, 	 -86, 	 -87, 	 -87, 	 -87, 	 -88, 	 -88, 	 -90, 	 -88, 	 -91, 	 -90, 	 -91, 	 -90, 	 -91, 	 -93, 	 -93, 	 -93, 	 -91, 	 -88, 	 -81, 	 -78, 	 -78, 	 -74, 	 -57, 	 -34, 	 -54, 	 -62, 	 -65, 	 -66, 	 -71, 	 -74, 	 -66, 	 -65, 	 -62, 	 -59, 	 -49, 	   5, 	  78, 	   4, 	 -27, 	 -30, 	 -32, 	 -35, 	 -35, 	 -32, 	 -34, 	 -35, 	 -37, 	 -40, 	 -42, 	 -66, 	 -65, 	 -68, 	 -71, 	 -71, 	 -59, 		  10, 	   3, 	 -57, 	 -75, 	 -77, 	 -74, 	 -69, 	 -71, 	 -70, 	 -60, 	 -60, 	  -9, 	  48, 	   5, 	 -82, 	 -86, 	 -85, 	 -86, 	 -89, 	 -88, 	 -87, 	 -88, 	 -86, 	 -90, 	 -90, 	 -91, 	 -89, 	 -88, 	 -73, 	 -51, 	 -11, 	 -20, 	 -72, 	 -49, 	  52, 	  54, 	  17, 	 -78, 	 -76, 	 -79, 	 -80, 	 -83, 	 -88, 	 -82, 	 -72, 	 -76, 	 -81, 	 -83, 	 -83, 	 -76, 	 -65, 	 -26, 	  41, 	  58, 	 -41, 	 -35, 	 -22, 	 -34, 	 -55, 	 -64, 	 -66, 	 -70, 	 -73, 	 -70, 	
 -65, 	 -73, 	 -81, 	 -83, 	 -84, 	 -85, 	 -85, 	 -84, 	 -85, 	 -87, 	 -86, 	 -87, 	 -87, 	 -88, 	 -87, 	 -88, 	 -88, 	 -90, 	 -90, 	 -91, 	 -93, 	 -92, 	 -93, 	 -93, 	 -92, 	 -91, 	 -90, 	 -88, 	 -79, 	 -77, 	 -79, 	 -73, 	 -48, 	 -35, 	 -57, 	 -63, 	 -64, 	 -67, 	 -72, 	 -67, 	 -67, 	 -65, 	 -62, 	 -52, 	 -27, 	  65, 	  39, 	 -26, 	 -31, 	 -34, 	 -38, 	 -30, 	 -36, 	 -33, 	 -37, 	 -38, 	 -37, 	 -40, 	 -62, 	 -68, 	 -66, 	 -70, 	 -69, 	 -63, 		 -18, 	  15, 	 -38, 	 -67, 	 -71, 	 -73, 	 -71, 	 -74, 	 -69, 	 -66, 	 -66, 	 -34, 	  37, 	  14, 	 -81, 	 -86, 	 -90, 	 -86, 	 -89, 	 -90, 	 -91, 	 -91, 	 -89, 	 -89, 	 -91, 	 -90, 	 -92, 	 -85, 	 -78, 	 -27, 	  20, 	 -52, 	 -65, 	 -35, 	  46, 	  50, 	  48, 	  -9, 	 -65, 	 -76, 	 -81, 	 -83, 	 -83, 	 -79, 	 -73, 	 -79, 	 -82, 	 -77, 	 -82, 	 -81, 	 -54, 	  15, 	  77, 	 -19, 	 -59, 	 -47, 	 -29, 	 -47, 	 -66, 	 -69, 	 -73, 	 -75, 	 -77, 	 -73, 	
 -48, 	 -61, 	 -72, 	 -78, 	 -84, 	 -80, 	 -84, 	 -81, 	 -84, 	 -85, 	 -86, 	 -84, 	 -85, 	 -81, 	 -86, 	 -89, 	 -89, 	 -90, 	 -90, 	 -90, 	 -91, 	 -92, 	 -91, 	 -94, 	 -93, 	 -93, 	 -92, 	 -92, 	 -86, 	 -79, 	 -79, 	 -76, 	 -69, 	 -37, 	 -42, 	 -61, 	 -64, 	 -68, 	 -71, 	 -67, 	 -66, 	 -67, 	 -64, 	 -58, 	 -40, 	  29, 	  73, 	 -10, 	 -29, 	 -33, 	 -33, 	 -32, 	 -34, 	 -41, 	 -30, 	 -37, 	 -39, 	 -41, 	 -47, 	 -68, 	 -68, 	 -72, 	 -71, 	 -70, 		 -46, 	  18, 	 -18, 	 -65, 	 -66, 	 -74, 	 -74, 	 -74, 	 -71, 	 -73, 	 -79, 	 -69, 	 -19, 	 -52, 	 -83, 	 -84, 	 -87, 	 -88, 	 -88, 	 -89, 	 -89, 	 -90, 	 -90, 	 -89, 	 -90, 	 -91, 	 -88, 	 -85, 	 -75, 	 -80, 	 -77, 	 -73, 	 -54, 	  21, 	  61, 	  61, 	  52, 	   0, 	 -58, 	 -78, 	 -81, 	 -84, 	 -82, 	 -77, 	 -76, 	 -83, 	 -82, 	 -77, 	 -81, 	 -74, 	 -57, 	  -4, 	  23, 	 -55, 	 -70, 	 -59, 	 -46, 	 -56, 	 -68, 	 -71, 	 -74, 	 -75, 	 -77, 	 -73, 	
 -25, 	 -26, 	 -39, 	 -65, 	 -77, 	 -77, 	 -78, 	 -82, 	 -80, 	 -82, 	 -83, 	 -83, 	 -78, 	 -77, 	 -80, 	 -87, 	 -88, 	 -89, 	 -89, 	 -90, 	 -91, 	 -91, 	 -92, 	 -93, 	 -93, 	 -92, 	 -92, 	 -92, 	 -90, 	 -83, 	 -79, 	 -78, 	 -76, 	 -64, 	 -29, 	 -52, 	 -63, 	 -65, 	 -68, 	 -69, 	 -67, 	 -63, 	 -65, 	 -62, 	 -46, 	 -15, 	  77, 	  25, 	 -26, 	 -32, 	 -33, 	 -35, 	 -35, 	 -34, 	 -38, 	 -36, 	 -37, 	 -40, 	 -48, 	 -65, 	 -71, 	 -73, 	 -73, 	 -71, 		 -63, 	   2, 	   0, 	 -53, 	 -73, 	 -69, 	 -74, 	 -73, 	 -72, 	 -76, 	 -85, 	 -84, 	 -83, 	 -84, 	 -88, 	 -88, 	 -87, 	 -87, 	 -88, 	 -90, 	 -90, 	 -89, 	 -90, 	 -89, 	 -90, 	 -89, 	 -86, 	 -82, 	 -80, 	 -79, 	 -77, 	 -60, 	  16, 	  45, 	  62, 	  58, 	  49, 	  34, 	 -64, 	 -79, 	 -82, 	 -81, 	 -81, 	 -74, 	 -76, 	 -86, 	 -83, 	 -77, 	 -78, 	 -74, 	 -60, 	 -44, 	 -50, 	 -55, 	 -69, 	 -69, 	 -67, 	 -64, 	 -70, 	 -76, 	 -78, 	 -75, 	 -72, 	 -71, 	
 -25, 	 -17, 	 -15, 	 -12, 	 -35, 	 -57, 	 -70, 	 -74, 	 -76, 	 -80, 	 -79, 	 -78, 	 -78, 	 -73, 	 -73, 	 -72, 	 -82, 	 -88, 	 -89, 	 -90, 	 -90, 	 -91, 	 -91, 	 -93, 	 -93, 	 -92, 	 -92, 	 -93, 	 -92, 	 -89, 	 -82, 	 -80, 	 -78, 	 -75, 	 -55, 	 -33, 	 -57, 	 -66, 	 -68, 	 -67, 	 -67, 	 -68, 	 -64, 	 -53, 	 -49, 	 -35, 	  51, 	  68, 	 -18, 	 -32, 	 -34, 	 -33, 	 -32, 	 -39, 	 -35, 	 -38, 	 -38, 	 -35, 	 -40, 	 -56, 	 -68, 	 -50, 	 -63, 	 -71, 		 -70, 	 -31, 	  17, 	 -33, 	 -69, 	 -73, 	 -70, 	 -71, 	 -80, 	 -77, 	 -77, 	 -77, 	 -81, 	 -86, 	 -85, 	 -87, 	 -88, 	 -87, 	 -89, 	 -89, 	 -89, 	 -88, 	 -88, 	 -89, 	 -90, 	 -87, 	 -82, 	 -83, 	 -81, 	 -82, 	 -71, 	 -52, 	  28, 	  40, 	  56, 	  64, 	  53, 	  50, 	 -39, 	 -77, 	 -80, 	 -80, 	 -81, 	 -73, 	 -80, 	 -85, 	 -85, 	 -81, 	 -81, 	 -73, 	 -66, 	 -50, 	 -64, 	 -62, 	 -64, 	 -73, 	 -71, 	 -68, 	 -71, 	 -77, 	 -78, 	 -73, 	 -71, 	 -72, 	
 -26, 	 -19, 	 -15, 	  -7, 	  -5, 	  -8, 	 -24, 	 -44, 	 -66, 	 -71, 	 -74, 	 -73, 	 -74, 	 -69, 	 -68, 	 -66, 	 -67, 	 -81, 	 -90, 	 -92, 	 -89, 	 -91, 	 -91, 	 -91, 	 -90, 	 -93, 	 -91, 	 -94, 	 -93, 	 -92, 	 -87, 	 -80, 	 -78, 	 -79, 	 -71, 	 -46, 	 -37, 	 -49, 	 -66, 	 -67, 	 -69, 	 -67, 	 -67, 	 -59, 	 -56, 	 -51, 	   8, 	  82, 	  15, 	 -23, 	 -31, 	 -27, 	 -31, 	 -34, 	 -33, 	 -35, 	 -38, 	 -27, 	 -42, 	 -47, 	 -70, 	 -45, 	 -56, 	 -69, 		 -71, 	 -54, 	   7, 	 -12, 	 -50, 	 -73, 	 -73, 	 -81, 	 -83, 	 -83, 	 -78, 	 -83, 	 -86, 	 -86, 	 -88, 	 -86, 	 -91, 	 -87, 	 -89, 	 -87, 	 -87, 	 -86, 	 -88, 	 -85, 	 -86, 	 -84, 	 -84, 	 -83, 	 -79, 	 -77, 	 -69, 	 -55, 	  25, 	  41, 	  53, 	  60, 	  59, 	  52, 	   4, 	 -77, 	 -80, 	 -80, 	 -80, 	 -74, 	 -74, 	 -88, 	 -84, 	 -82, 	 -79, 	 -71, 	 -63, 	 -44, 	 -57, 	 -65, 	 -66, 	 -72, 	 -76, 	 -74, 	 -75, 	 -78, 	 -76, 	 -72, 	 -71, 	 -72, 	
 -33, 	 -29, 	 -18, 	  -9, 	  -8, 	  -2, 	  -7, 	 -13, 	 -23, 	 -42, 	 -63, 	 -66, 	 -68, 	 -66, 	 -62, 	 -65, 	 -66, 	 -71, 	 -83, 	 -89, 	 -91, 	 -88, 	 -90, 	 -90, 	 -92, 	 -91, 	 -92, 	 -91, 	 -92, 	 -91, 	 -91, 	 -87, 	 -80, 	 -77, 	 -77, 	 -67, 	 -33, 	 -45, 	 -56, 	 -65, 	 -69, 	 -64, 	 -67, 	 -62, 	 -61, 	 -59, 	 -22, 	  66, 	  57, 	 -21, 	 -29, 	 -26, 	 -27, 	 -31, 	 -38, 	 -36, 	 -35, 	 -35, 	 -34, 	 -39, 	 -65, 	 -66, 	 -62, 	 -68, 		 -71, 	 -63, 	 -19, 	 -12, 	 -50, 	 -76, 	 -82, 	 -79, 	 -82, 	 -81, 	 -84, 	 -86, 	 -81, 	 -81, 	 -83, 	 -82, 	 -80, 	 -81, 	 -83, 	 -80, 	 -77, 	 -75, 	 -76, 	 -77, 	 -77, 	 -76, 	 -76, 	 -75, 	 -74, 	 -70, 	 -66, 	 -57, 	  12, 	  44, 	  48, 	  58, 	  63, 	  53, 	  34, 	 -65, 	 -79, 	 -79, 	 -76, 	 -64, 	 -77, 	 -86, 	 -83, 	 -83, 	 -80, 	 -71, 	 -65, 	 -49, 	 -61, 	 -64, 	 -71, 	 -75, 	 -78, 	 -77, 	 -78, 	 -78, 	 -75, 	 -70, 	 -70, 	 -73, 	
 -32, 	 -29, 	 -26, 	 -19, 	 -12, 	 -11, 	  -6, 	  -7, 	 -12, 	 -21, 	 -34, 	 -51, 	 -60, 	 -61, 	 -60, 	 -60, 	 -62, 	 -66, 	 -78, 	 -86, 	 -90, 	 -90, 	 -90, 	 -89, 	 -91, 	 -91, 	 -91, 	 -92, 	 -93, 	 -91, 	 -91, 	 -89, 	 -84, 	 -79, 	 -77, 	 -76, 	 -58, 	 -30, 	 -55, 	 -64, 	 -67, 	 -64, 	 -64, 	 -60, 	 -64, 	 -63, 	 -44, 	  25, 	  84, 	   4, 	 -25, 	 -27, 	 -28, 	 -36, 	 -36, 	 -37, 	 -35, 	 -34, 	 -31, 	 -44, 	 -53, 	 -67, 	 -43, 	 -64, 		 -68, 	 -69, 	 -52, 	 -33, 	 -67, 	 -76, 	 -77, 	 -78, 	 -81, 	 -77, 	 -71, 	 -70, 	 -30, 	 -54, 	 -68, 	 -69, 	 -68, 	 -69, 	 -70, 	 -68, 	 -68, 	 -65, 	 -65, 	 -65, 	 -63, 	 -67, 	 -65, 	 -66, 	 -66, 	 -67, 	 -63, 	 -59, 	   4, 	  40, 	  46, 	  52, 	  65, 	  56, 	  49, 	 -24, 	 -79, 	 -80, 	 -73, 	 -67, 	 -75, 	 -87, 	 -87, 	 -85, 	 -75, 	 -70, 	 -66, 	 -50, 	 -61, 	 -69, 	 -69, 	 -76, 	 -79, 	 -81, 	 -81, 	 -76, 	 -70, 	 -69, 	 -68, 	 -73, 	
 -39, 	 -31, 	 -29, 	 -22, 	 -19, 	 -15, 	 -13, 	  -8, 	 -14, 	 -19, 	 -30, 	 -40, 	 -43, 	 -54, 	 -53, 	 -58, 	 -62, 	 -68, 	 -72, 	 -79, 	 -85, 	 -88, 	 -87, 	 -88, 	 -88, 	 -87, 	 -92, 	 -90, 	 -92, 	 -92, 	 -90, 	 -91, 	 -88, 	 -81, 	 -79, 	 -80, 	 -76, 	 -50, 	 -34, 	 -63, 	 -66, 	 -63, 	 -62, 	 -62, 	 -67, 	 -65, 	 -50, 	  -7, 	  90, 	  40, 	 -24, 	 -31, 	 -30, 	 -34, 	 -38, 	 -37, 	 -35, 	 -29, 	 -36, 	 -44, 	 -48, 	 -58, 	 -56, 	 -45, 		 -52, 	 -64, 	 -65, 	 -63, 	 -62, 	 -65, 	 -59, 	 -65, 	 -71, 	 -72, 	 -68, 	 -53, 	  35, 	  25, 	 -48, 	 -48, 	 -48, 	 -45, 	 -44, 	 -41, 	 -34, 	 -30, 	 -22, 	  -9, 	  -4, 	   4, 	 -21, 	 -29, 	 -32, 	 -46, 	 -43, 	 -45, 	  -4, 	  39, 	  41, 	  44, 	  59, 	  54, 	  51, 	  23, 	 -70, 	 -77, 	 -76, 	 -72, 	 -76, 	 -86, 	 -85, 	 -81, 	 -74, 	 -70, 	 -65, 	 -51, 	 -61, 	 -65, 	 -70, 	 -76, 	 -78, 	 -81, 	 -82, 	 -77, 	 -67, 	 -70, 	 -69, 	 -72, 	
 -31, 	 -32, 	 -34, 	 -29, 	 -20, 	 -13, 	 -17, 	 -19, 	 -19, 	 -24, 	 -29, 	 -40, 	 -44, 	 -48, 	 -52, 	 -52, 	 -56, 	 -65, 	 -72, 	 -78, 	 -84, 	 -86, 	 -87, 	 -87, 	 -87, 	 -89, 	 -88, 	 -90, 	 -91, 	 -90, 	 -90, 	 -91, 	 -90, 	 -85, 	 -80, 	 -78, 	 -76, 	 -69, 	 -33, 	 -44, 	 -62, 	 -65, 	 -64, 	 -64, 	 -67, 	 -66, 	 -47, 	 -28, 	  43, 	  76, 	 -15, 	 -30, 	 -30, 	 -33, 	 -35, 	 -34, 	 -36, 	 -35, 	 -35, 	 -38, 	 -46, 	 -55, 	 -64, 	 -60, 		 -14, 	 -40, 	 -68, 	 -71, 	 -63, 	   2, 	   9, 	 -50, 	 -61, 	 -63, 	 -57, 	 -47, 	  43, 	  58, 	  47, 	  42, 	  48, 	  47, 	  51, 	  48, 	  52, 	  57, 	  58, 	  60, 	  59, 	  58, 	  55, 	  55, 	  53, 	  40, 	  31, 	  18, 	   7, 	  37, 	  34, 	  32, 	  33, 	  45, 	  50, 	  49, 	 -48, 	 -78, 	 -71, 	 -72, 	 -78, 	 -82, 	 -88, 	 -80, 	 -71, 	 -64, 	 -67, 	 -45, 	 -54, 	 -63, 	 -73, 	 -78, 	 -80, 	 -81, 	 -82, 	 -78, 	 -70, 	 -69, 	 -70, 	 -73, 	
 -20, 	 -27, 	 -29, 	 -25, 	 -23, 	 -17, 	 -18, 	 -19, 	 -24, 	 -26, 	 -31, 	 -39, 	 -46, 	 -49, 	 -54, 	 -52, 	 -50, 	 -57, 	 -70, 	 -79, 	 -84, 	 -86, 	 -85, 	 -87, 	 -88, 	 -86, 	 -88, 	 -90, 	 -90, 	 -91, 	 -90, 	 -90, 	 -91, 	 -87, 	 -85, 	 -78, 	 -79, 	 -75, 	 -64, 	 -29, 	 -52, 	 -61, 	 -61, 	 -61, 	 -66, 	 -63, 	 -56, 	 -39, 	   1, 	  83, 	   8, 	 -21, 	 -33, 	 -31, 	 -37, 	 -33, 	 -33, 	 -30, 	 -31, 	 -36, 	 -42, 	 -45, 	 -59, 	 -70, 		 -68, 	 -55, 	 -72, 	 -72, 	 -62, 	 -15, 	  72, 	  38, 	 -17, 	   8, 	  -8, 	   9, 	  58, 	  67, 	  65, 	  63, 	  64, 	  62, 	  62, 	  61, 	  60, 	  61, 	  63, 	  63, 	  60, 	  56, 	  29, 	  21, 	  13, 	   7, 	  -6, 	   8, 	   1, 	   0, 	  -3, 	  -9, 	  -9, 	   8, 	  36, 	  48, 	  -1, 	 -72, 	 -70, 	 -71, 	 -75, 	 -82, 	 -83, 	 -74, 	 -69, 	 -64, 	 -66, 	 -47, 	 -55, 	 -62, 	 -73, 	 -77, 	 -81, 	 -79, 	 -81, 	 -79, 	 -73, 	 -70, 	 -68, 	 -71, 	
 -12, 	 -13, 	 -22, 	 -17, 	 -24, 	 -19, 	 -22, 	 -18, 	 -22, 	 -28, 	 -29, 	 -41, 	 -47, 	 -51, 	 -54, 	 -51, 	 -52, 	 -51, 	 -55, 	 -71, 	 -81, 	 -83, 	 -85, 	 -83, 	 -87, 	 -87, 	 -89, 	 -89, 	 -90, 	 -90, 	 -91, 	 -90, 	 -88, 	 -90, 	 -90, 	 -82, 	 -79, 	 -78, 	 -72, 	 -51, 	 -33, 	 -53, 	 -60, 	 -64, 	 -62, 	 -62, 	 -59, 	 -54, 	 -22, 	  63, 	  45, 	 -13, 	 -24, 	 -34, 	 -32, 	 -34, 	 -32, 	 -36, 	 -36, 	 -35, 	 -37, 	 -44, 	 -53, 	 -66, 		 -69, 	 -75, 	 -78, 	 -72, 	 -68, 	 -47, 	  30, 	  78, 	  70, 	  42, 	  28, 	  57, 	  64, 	  64, 	  66, 	  64, 	  64, 	  65, 	  66, 	  67, 	  61, 	  66, 	  68, 	  69, 	  67, 	  66, 	  58, 	  42, 	  50, 	  31, 	  13, 	 -13, 	  -9, 	 -20, 	 -21, 	 -25, 	 -19, 	   4, 	  31, 	  41, 	  27, 	 -57, 	 -62, 	 -71, 	 -77, 	 -78, 	 -83, 	 -71, 	 -63, 	 -68, 	 -66, 	 -53, 	 -58, 	 -70, 	 -72, 	 -78, 	 -80, 	 -78, 	 -77, 	 -77, 	 -76, 	 -71, 	 -69, 	 -72, 	
 -23, 	 -13, 	  -6, 	 -15, 	 -17, 	 -16, 	 -23, 	 -22, 	 -24, 	 -29, 	 -35, 	 -39, 	 -41, 	 -50, 	 -49, 	 -51, 	 -49, 	 -44, 	 -39, 	 -54, 	 -76, 	 -81, 	 -82, 	 -84, 	 -85, 	 -84, 	 -88, 	 -89, 	 -89, 	 -89, 	 -89, 	 -90, 	 -89, 	 -89, 	 -90, 	 -89, 	 -80, 	 -79, 	 -78, 	 -71, 	 -37, 	 -40, 	 -56, 	 -60, 	 -60, 	 -63, 	 -60, 	 -58, 	 -42, 	  20, 	  68, 	   6, 	 -23, 	 -25, 	 -30, 	 -36, 	 -34, 	 -32, 	 -37, 	 -37, 	 -31, 	 -36, 	 -46, 	 -64, 		 -66, 	 -70, 	 -76, 	 -74, 	 -71, 	 -61, 	 -24, 	  79, 	  81, 	  49, 	  12, 	  65, 	  73, 	  77, 	  77, 	  73, 	  69, 	  69, 	  69, 	  70, 	  69, 	  64, 	  71, 	  70, 	  75, 	  74, 	  68, 	  59, 	  56, 	  72, 	  65, 	  32, 	  -1, 	 -17, 	 -21, 	 -24, 	 -32, 	 -14, 	  40, 	  35, 	  33, 	 -18, 	 -67, 	 -73, 	 -74, 	 -79, 	 -82, 	 -75, 	 -64, 	 -63, 	 -66, 	 -54, 	 -63, 	 -72, 	 -75, 	 -78, 	 -78, 	 -75, 	 -72, 	 -77, 	 -74, 	 -76, 	 -74, 	 -73, 	
 -42, 	 -39, 	 -29, 	 -16, 	 -13, 	 -18, 	 -22, 	 -19, 	 -28, 	 -29, 	 -31, 	 -35, 	 -39, 	 -46, 	 -50, 	 -48, 	 -46, 	 -44, 	 -39, 	 -32, 	 -51, 	 -78, 	 -80, 	 -83, 	 -82, 	 -85, 	 -85, 	 -87, 	 -88, 	 -89, 	 -88, 	 -89, 	 -88, 	 -89, 	 -89, 	 -89, 	 -86, 	 -81, 	 -77, 	 -76, 	 -67, 	 -32, 	 -51, 	 -58, 	 -59, 	 -61, 	 -62, 	 -54, 	 -50, 	 -27, 	  68, 	  32, 	 -22, 	 -30, 	 -28, 	 -31, 	 -32, 	 -34, 	 -32, 	 -37, 	 -28, 	 -28, 	 -39, 	 -58, 		 -64, 	 -66, 	 -73, 	 -76, 	 -74, 	 -71, 	 -56, 	  23, 	  81, 	  63, 	   9, 	  47, 	  78, 	  78, 	  79, 	  77, 	  72, 	  73, 	  73, 	  67, 	  70, 	  67, 	  67, 	  71, 	  76, 	  75, 	  74, 	  71, 	  68, 	  74, 	  75, 	  46, 	   3, 	  -9, 	 -14, 	 -15, 	 -28, 	 -22, 	  36, 	  39, 	  42, 	   3, 	 -65, 	 -73, 	 -73, 	 -78, 	 -83, 	 -71, 	 -61, 	 -58, 	 -66, 	 -58, 	 -61, 	 -71, 	 -79, 	 -77, 	 -73, 	 -70, 	 -72, 	 -76, 	 -74, 	 -76, 	 -77, 	 -75, 	

 -59, 	 -53, 	 -50, 	 -43, 	 -33, 	 -17, 	 -19, 	 -23, 	 -29, 	 -30, 	 -34, 	 -39, 	 -37, 	 -42, 	 -45, 	 -48, 	 -44, 	 -41, 	 -36, 	 -35, 	 -26, 	 -51, 	 -79, 	 -78, 	 -81, 	 -82, 	 -84, 	 -85, 	 -85, 	 -87, 	 -86, 	 -87, 	 -87, 	 -87, 	 -89, 	 -90, 	 -87, 	 -82, 	 -80, 	 -75, 	 -74, 	 -56, 	 -35, 	 -53, 	 -47, 	 -60, 	 -60, 	 -59, 	 -57, 	 -41, 	  33, 	  69, 	 -14, 	 -29, 	 -22, 	 -31, 	 -34, 	 -29, 	 -34, 	 -32, 	 -33, 	 -32, 	 -38, 	 -49, 		 -61, 	 -64, 	 -73, 	 -68, 	 -70, 	 -73, 	 -64, 	 -43, 	  58, 	  74, 	  26, 	  14, 	  54, 	  47, 	  51, 	  66, 	  75, 	  73, 	  70, 	  62, 	  63, 	  74, 	  68, 	  72, 	  63, 	  74, 	  74, 	  72, 	  76, 	  75, 	  72, 	  62, 	  11, 	  12, 	 -10, 	 -16, 	 -17, 	 -23, 	  10, 	  37, 	  40, 	  34, 	 -49, 	 -72, 	 -73, 	 -78, 	 -79, 	 -68, 	 -55, 	 -57, 	 -62, 	 -54, 	 -58, 	 -69, 	 -60, 	 -32, 	 -10, 	 -25, 	 -49, 	 -58, 	 -74, 	 -76, 	 -72, 	 -79, 	
 -62, 	 -62, 	 -62, 	 -57, 	 -50, 	 -40, 	 -29, 	 -27, 	 -29, 	 -36, 	 -40, 	 -43, 	 -38, 	 -40, 	 -42, 	 -46, 	 -44, 	 -41, 	 -36, 	 -28, 	 -24, 	 -23, 	 -53, 	 -77, 	 -79, 	 -83, 	 -83, 	 -84, 	 -85, 	 -86, 	 -85, 	 -87, 	 -87, 	 -87, 	 -90, 	 -90, 	 -88, 	 -89, 	 -83, 	 -78, 	 -79, 	 -72, 	 -39, 	 -41, 	 -48, 	 -59, 	 -57, 	 -62, 	 -59, 	 -51, 	  -3, 	  74, 	  15, 	 -27, 	 -31, 	 -26, 	 -33, 	 -31, 	 -33, 	 -33, 	 -31, 	 -33, 	 -39, 	 -43, 		 -57, 	 -61, 	 -67, 	 -52, 	 -42, 	 -65, 	 -69, 	 -67, 	 -17, 	  77, 	  29, 	  -7, 	  25, 	  -1, 	  32, 	  57, 	  71, 	  74, 	  47, 	  60, 	  31, 	  63, 	  67, 	  68, 	  56, 	  58, 	  71, 	  72, 	  72, 	  69, 	  74, 	  68, 	  41, 	  24, 	   3, 	 -17, 	 -17, 	 -18, 	 -10, 	  24, 	  35, 	  36, 	 -18, 	 -71, 	 -72, 	 -77, 	 -77, 	 -64, 	 -53, 	 -63, 	 -69, 	 -55, 	 -56, 	 -70, 	 -64, 	 -25, 	  -1, 	  18, 	   6, 	 -45, 	 -55, 	 -73, 	 -72, 	 -76, 	
 -55, 	 -60, 	 -60, 	 -61, 	 -58, 	 -50, 	 -43, 	 -37, 	 -31, 	 -37, 	 -40, 	 -41, 	 -44, 	 -46, 	 -43, 	 -41, 	 -42, 	 -39, 	 -33, 	 -25, 	 -21, 	 -17, 	 -21, 	 -48, 	 -75, 	 -79, 	 -81, 	 -83, 	 -81, 	 -82, 	 -83, 	 -86, 	 -86, 	 -86, 	 -89, 	 -89, 	 -92, 	 -87, 	 -85, 	 -80, 	 -81, 	 -78, 	 -63, 	 -31, 	 -46, 	 -55, 	 -58, 	 -60, 	 -61, 	 -57, 	 -32, 	  48, 	  39, 	 -16, 	 -28, 	 -26, 	 -31, 	 -26, 	 -34, 	 -30, 	 -34, 	 -29, 	 -39, 	 -41, 		 -52, 	 -57, 	 -61, 	 -48, 	 -28, 	 -46, 	 -69, 	 -73, 	 -64, 	 -18, 	 -12, 	 -22, 	  -6, 	 -21, 	  10, 	  58, 	  63, 	  64, 	  57, 	  60, 	  50, 	  59, 	  65, 	  65, 	  66, 	  54, 	  58, 	  60, 	  57, 	  54, 	  64, 	  70, 	  55, 	  22, 	   9, 	 -14, 	  -8, 	 -10, 	  -7, 	  15, 	  36, 	  38, 	  20, 	 -68, 	 -70, 	 -80, 	 -72, 	 -61, 	 -62, 	 -70, 	 -69, 	 -58, 	 -65, 	 -83, 	 -78, 	 -59, 	 -31, 	 -32, 	 -19, 	 -41, 	 -53, 	 -66, 	 -72, 	 -77, 	
 -51, 	 -55, 	 -56, 	 -57, 	 -56, 	 -57, 	 -57, 	 -46, 	 -41, 	 -40, 	 -44, 	 -41, 	 -44, 	 -44, 	 -42, 	 -43, 	 -40, 	 -38, 	 -32, 	 -23, 	 -18, 	 -12, 	 -16, 	 -18, 	 -51, 	 -74, 	 -81, 	 -79, 	 -75, 	 -71, 	 -77, 	 -81, 	 -86, 	 -85, 	 -88, 	 -89, 	 -88, 	 -90, 	 -89, 	 -81, 	 -78, 	 -78, 	 -75, 	 -48, 	 -32, 	 -54, 	 -56, 	 -60, 	 -63, 	 -58, 	 -38, 	   9, 	  67, 	   2, 	 -22, 	 -24, 	 -27, 	 -28, 	 -27, 	 -30, 	 -29, 	 -30, 	 -34, 	 -42, 		 -46, 	 -57, 	 -56, 	 -49, 	 -28, 	 -45, 	 -64, 	 -72, 	 -72, 	 -63, 	 -35, 	 -22, 	 -24, 	 -25, 	 -14, 	  23, 	  62, 	  55, 	  54, 	  59, 	  69, 	  65, 	  63, 	  58, 	  65, 	  62, 	  57, 	  51, 	  54, 	  42, 	  48, 	  66, 	  59, 	  25, 	   8, 	 -10, 	 -15, 	  -7, 	   8, 	   7, 	  31, 	  39, 	  36, 	 -38, 	 -73, 	 -80, 	 -72, 	 -65, 	 -66, 	 -69, 	 -76, 	 -68, 	 -42, 	 -40, 	 -62, 	 -66, 	 -48, 	 -43, 	 -34, 	 -46, 	 -59, 	 -67, 	 -74, 	 -73, 	
 -54, 	 -51, 	 -52, 	 -51, 	 -52, 	 -52, 	 -52, 	 -54, 	 -52, 	 -41, 	 -41, 	 -47, 	 -46, 	 -40, 	 -39, 	 -38, 	 -35, 	 -33, 	 -28, 	 -22, 	 -16, 	 -14, 	 -10, 	 -15, 	 -19, 	 -57, 	 -70, 	 -75, 	 -73, 	 -68, 	 -65, 	 -77, 	 -81, 	 -86, 	 -88, 	 -88, 	 -92, 	 -91, 	 -91, 	 -87, 	 -82, 	 -79, 	 -76, 	 -69, 	 -38, 	 -41, 	 -55, 	 -62, 	 -60, 	 -58, 	 -49, 	 -16, 	  66, 	  30, 	 -21, 	 -25, 	 -25, 	 -26, 	 -27, 	 -26, 	 -31, 	 -33, 	 -35, 	 -39, 		 -41, 	 -52, 	 -58, 	 -45, 	 -23, 	 -42, 	 -55, 	 -60, 	 -63, 	 -56, 	 -47, 	 -27, 	 -29, 	 -31, 	 -36, 	  -8, 	  52, 	  62, 	  53, 	  61, 	  68, 	  66, 	  64, 	  54, 	  62, 	  61, 	  49, 	  46, 	  56, 	  50, 	  45, 	  61, 	  63, 	  35, 	   8, 	   3, 	   0, 	  -7, 	   2, 	   5, 	  25, 	  36, 	  38, 	  -2, 	 -72, 	 -75, 	 -65, 	 -62, 	 -65, 	 -71, 	 -73, 	 -76, 	 -73, 	 -55, 	 -64, 	 -67, 	 -56, 	 -51, 	 -43, 	 -54, 	 -66, 	 -68, 	 -70, 	 -74, 	
 -56, 	 -52, 	 -52, 	 -50, 	 -50, 	 -50, 	 -51, 	 -48, 	 -55, 	 -52, 	 -49, 	 -41, 	 -47, 	 -42, 	 -37, 	 -31, 	 -29, 	 -28, 	 -22, 	 -21, 	 -16, 	 -11, 	  -9, 	 -12, 	 -12, 	 -22, 	 -52, 	 -66, 	 -72, 	 -65, 	 -63, 	 -61, 	 -78, 	 -81, 	 -87, 	 -89, 	 -89, 	 -91, 	 -91, 	 -91, 	 -86, 	 -77, 	 -79, 	 -76, 	 -59, 	 -32, 	 -56, 	 -62, 	 -61, 	 -56, 	 -48, 	 -31, 	  36, 	  71, 	 -16, 	 -26, 	 -24, 	 -28, 	 -27, 	 -24, 	 -32, 	 -34, 	 -34, 	 -39, 		 -36, 	 -45, 	 -60, 	 -54, 	 -40, 	 -45, 	 -53, 	 -55, 	 -55, 	 -55, 	 -41, 	 -22, 	 -35, 	 -31, 	 -38, 	 -22, 	  20, 	  59, 	  54, 	  63, 	  63, 	  67, 	  66, 	  57, 	  56, 	  61, 	  48, 	  44, 	  55, 	  55, 	  45, 	  56, 	  63, 	  47, 	  32, 	  12, 	   6, 	   2, 	   8, 	   5, 	  13, 	  29, 	  32, 	  25, 	 -54, 	 -74, 	 -67, 	 -63, 	 -71, 	 -74, 	 -76, 	 -75, 	 -78, 	 -85, 	 -85, 	 -68, 	 -64, 	 -73, 	 -70, 	 -73, 	 -77, 	 -76, 	 -72, 	 -76, 	
 -56, 	 -57, 	 -52, 	 -52, 	 -47, 	 -46, 	 -44, 	 -47, 	 -47, 	 -53, 	 -55, 	 -51, 	 -47, 	 -45, 	 -39, 	 -27, 	 -15, 	 -15, 	 -16, 	 -13, 	 -12, 	 -13, 	  -6, 	  -9, 	  -8, 	 -17, 	 -32, 	 -60, 	 -61, 	 -65, 	 -61, 	 -59, 	 -64, 	 -83, 	 -85, 	 -88, 	 -88, 	 -91, 	 -91, 	 -90, 	 -90, 	 -84, 	 -81, 	 -78, 	 -73, 	 -49, 	 -37, 	 -59, 	 -55, 	 -57, 	 -49, 	 -44, 	   6, 	  84, 	  17, 	 -22, 	 -27, 	 -33, 	 -28, 	 -28, 	 -31, 	 -35, 	 -36, 	 -36, 		 -37, 	 -39, 	 -56, 	 -58, 	 -54, 	 -50, 	 -53, 	 -52, 	 -51, 	 -50, 	 -48, 	 -42, 	 -43, 	 -35, 	 -28, 	 -26, 	  -7, 	  46, 	  55, 	  51, 	  54, 	  61, 	  60, 	  56, 	  55, 	  54, 	  51, 	  42, 	  40, 	  43, 	  43, 	  55, 	  64, 	  50, 	  40, 	  18, 	   9, 	   8, 	  10, 	  11, 	   5, 	  23, 	  36, 	  34, 	 -11, 	 -68, 	 -68, 	 -71, 	 -74, 	 -73, 	 -77, 	 -78, 	 -82, 	 -80, 	 -74, 	 -72, 	 -79, 	 -84, 	 -86, 	 -83, 	 -79, 	 -75, 	 -76, 	 -76, 	
 -56, 	 -56, 	 -55, 	 -50, 	 -48, 	 -45, 	 -39, 	 -39, 	 -42, 	 -46, 	 -48, 	 -53, 	 -55, 	 -52, 	 -44, 	 -38, 	 -20, 	  -7, 	  -8, 	  -8, 	  -7, 	  -7, 	  -8, 	  -7, 	 -10, 	 -17, 	 -22, 	 -39, 	 -52, 	 -55, 	 -58, 	 -53, 	 -56, 	 -72, 	 -87, 	 -87, 	 -91, 	 -90, 	 -91, 	 -91, 	 -92, 	 -89, 	 -81, 	 -78, 	 -78, 	 -68, 	 -34, 	 -52, 	 -57, 	 -56, 	 -53, 	 -47, 	 -27, 	  60, 	  60, 	 -19, 	 -29, 	 -34, 	 -32, 	 -30, 	 -34, 	 -28, 	 -32, 	 -34, 		 -42, 	 -46, 	 -51, 	 -58, 	 -55, 	 -52, 	 -52, 	 -49, 	 -49, 	 -53, 	 -51, 	 -46, 	 -46, 	 -32, 	 -17, 	 -12, 	  -1, 	   4, 	  44, 	  57, 	  43, 	  37, 	  65, 	  53, 	  46, 	  45, 	  51, 	  25, 	  26, 	  11, 	  21, 	  49, 	  64, 	  50, 	  44, 	  29, 	   9, 	   5, 	  11, 	  14, 	  19, 	  19, 	  37, 	  38, 	  27, 	 -27, 	 -65, 	 -70, 	 -74, 	 -78, 	 -78, 	 -75, 	 -75, 	 -80, 	 -82, 	 -85, 	 -87, 	 -83, 	 -75, 	 -71, 	 -71, 	 -75, 	 -73, 	 -75, 	
 -55, 	 -59, 	 -52, 	 -52, 	 -49, 	 -47, 	 -44, 	 -35, 	 -36, 	 -37, 	 -47, 	 -51, 	 -52, 	 -58, 	 -57, 	 -45, 	 -35, 	 -16, 	  -4, 	   0, 	  -1, 	  -6, 	  -8, 	 -13, 	  -9, 	 -16, 	 -22, 	 -32, 	 -42, 	 -48, 	 -48, 	 -53, 	 -54, 	 -61, 	 -84, 	 -89, 	 -88, 	 -91, 	 -90, 	 -91, 	 -90, 	 -90, 	 -84, 	 -78, 	 -79, 	 -72, 	 -55, 	 -32, 	 -59, 	 -58, 	 -54, 	 -54, 	 -41, 	  20, 	  93, 	   3, 	 -27, 	 -34, 	 -35, 	 -33, 	 -29, 	 -26, 	 -30, 	 -27, 		 -37, 	 -42, 	 -50, 	 -60, 	 -62, 	 -59, 	 -51, 	 -53, 	 -51, 	 -50, 	 -48, 	 -44, 	 -45, 	 -34, 	 -13, 	 -15, 	 -17, 	 -17, 	 -20, 	  31, 	  55, 	  35, 	  69, 	  53, 	  41, 	  40, 	  52, 	  25, 	  18, 	   8, 	  19, 	  37, 	  56, 	  59, 	  52, 	  44, 	  22, 	  14, 	  16, 	   5, 	   9, 	  30, 	  35, 	  40, 	  35, 	 -14, 	 -53, 	 -65, 	 -73, 	 -79, 	 -79, 	 -74, 	 -71, 	 -71, 	 -76, 	 -81, 	 -81, 	 -73, 	 -67, 	 -68, 	 -70, 	 -73, 	 -73, 	 -74, 	
 -58, 	 -62, 	 -59, 	 -53, 	 -49, 	 -50, 	 -45, 	 -40, 	 -34, 	 -36, 	 -42, 	 -49, 	 -50, 	 -53, 	 -60, 	 -59, 	 -47, 	 -37, 	 -19, 	  -3, 	   0, 	  -5, 	  -8, 	 -15, 	 -14, 	 -18, 	 -23, 	 -31, 	 -36, 	 -39, 	 -42, 	 -47, 	 -55, 	 -65, 	 -76, 	 -88, 	 -90, 	 -90, 	 -89, 	 -90, 	 -91, 	 -92, 	 -90, 	 -81, 	 -80, 	 -78, 	 -65, 	 -40, 	 -44, 	 -48, 	 -46, 	 -41, 	 -41, 	  -6, 	  97, 	  50, 	 -24, 	 -34, 	 -39, 	 -33, 	 -30, 	 -33, 	 -24, 	 -27, 		 -27, 	 -38, 	 -40, 	 -55, 	 -63, 	 -67, 	 -62, 	 -57, 	 -49, 	 -49, 	 -43, 	 -32, 	 -42, 	 -37, 	 -25, 	 -14, 	 -35, 	 -31, 	 -31, 	   3, 	  57, 	  49, 	  56, 	  47, 	  46, 	  33, 	  45, 	  33, 	  23, 	  16, 	  19, 	  29, 	  55, 	  62, 	  58, 	  48, 	  28, 	  18, 	  15, 	   2, 	   4, 	  28, 	  39, 	  39, 	  33, 	   4, 	 -54, 	 -68, 	 -73, 	 -74, 	 -73, 	 -71, 	 -69, 	 -66, 	 -62, 	 -65, 	 -61, 	 -59, 	 -61, 	 -64, 	 -68, 	 -73, 	 -68, 	 -67, 	
 -59, 	 -61, 	 -61, 	 -57, 	 -53, 	 -49, 	 -47, 	 -44, 	 -40, 	 -34, 	 -34, 	 -42, 	 -48, 	 -54, 	 -52, 	 -61, 	 -58, 	 -52, 	 -38, 	 -22, 	  -4, 	  -3, 	 -14, 	 -15, 	 -16, 	 -20, 	 -23, 	 -30, 	 -29, 	 -40, 	 -43, 	 -47, 	 -55, 	 -69, 	 -76, 	 -84, 	 -89, 	 -89, 	 -89, 	 -89, 	 -91, 	 -91, 	 -90, 	 -85, 	 -81, 	 -81, 	 -76, 	 -64, 	 -27, 	 -35, 	 -48, 	 -53, 	 -42, 	 -28, 	  65, 	  83, 	 -18, 	 -26, 	 -33, 	 -36, 	 -34, 	 -30, 	 -32, 	 -25, 		 -27, 	 -38, 	 -40, 	 -42, 	 -63, 	 -65, 	 -61, 	 -56, 	 -51, 	 -50, 	 -47, 	 -29, 	 -29, 	 -36, 	 -29, 	 -16, 	 -17, 	 -27, 	  -2, 	   9, 	  46, 	  60, 	  55, 	  41, 	  33, 	  44, 	  48, 	  48, 	  42, 	  39, 	  28, 	  35, 	  47, 	  60, 	  58, 	  49, 	  33, 	  25, 	  18, 	   7, 	  -4, 	  10, 	  42, 	  36, 	  38, 	  24, 	 -50, 	 -69, 	 -72, 	 -72, 	 -67, 	 -65, 	 -60, 	 -58, 	 -52, 	 -57, 	 -54, 	 -43, 	 -44, 	 -49, 	 -46, 	 -39, 	 -26, 	 -18, 	
 -61, 	 -61, 	 -59, 	 -59, 	 -58, 	 -55, 	 -52, 	 -47, 	 -42, 	 -36, 	 -39, 	 -39, 	 -42, 	 -50, 	 -50, 	 -54, 	 -60, 	 -60, 	 -53, 	 -39, 	 -28, 	  -9, 	 -13, 	 -21, 	 -22, 	 -24, 	 -26, 	 -32, 	 -35, 	 -41, 	 -47, 	 -51, 	 -55, 	 -67, 	 -74, 	 -83, 	 -88, 	 -87, 	 -90, 	 -89, 	 -90, 	 -91, 	 -90, 	 -89, 	 -82, 	 -77, 	 -78, 	 -75, 	 -38, 	 -32, 	 -56, 	 -59, 	 -49, 	 -42, 	  12, 	  95, 	  12, 	 -26, 	 -30, 	 -33, 	 -37, 	 -30, 	 -30, 	 -25, 		 -25, 	 -34, 	 -35, 	 -33, 	 -51, 	 -58, 	 -58, 	 -58, 	 -53, 	 -51, 	 -46, 	 -38, 	 -28, 	 -29, 	 -28, 	 -18, 	   2, 	  11, 	  17, 	  20, 	  42, 	  60, 	  59, 	  62, 	  62, 	  62, 	  57, 	  62, 	  52, 	  51, 	  44, 	  42, 	  45, 	  57, 	  59, 	  48, 	  42, 	  24, 	  29, 	  12, 	   0, 	   5, 	  41, 	  44, 	  48, 	  32, 	 -23, 	 -65, 	 -59, 	 -39, 	 -20, 	 -10, 	  -6, 	  -5, 	  -5, 	  -1, 	   9, 	  -1, 	  -2, 	  -8, 	  -7, 	 -13, 	 -26, 	 -33, 	
 -65, 	 -60, 	 -57, 	 -63, 	 -61, 	 -57, 	 -61, 	 -53, 	 -50, 	 -42, 	 -36, 	 -38, 	 -39, 	 -42, 	 -46, 	 -48, 	 -51, 	 -57, 	 -60, 	 -52, 	 -46, 	 -32, 	 -21, 	 -25, 	 -28, 	 -28, 	 -31, 	 -33, 	 -36, 	 -42, 	 -48, 	 -49, 	 -54, 	 -64, 	 -76, 	 -81, 	 -85, 	 -86, 	 -90, 	 -88, 	 -89, 	 -89, 	 -90, 	 -91, 	 -87, 	 -78, 	 -76, 	 -77, 	 -63, 	 -26, 	 -49, 	 -54, 	 -55, 	 -44, 	 -24, 	  63, 	  34, 	 -22, 	 -24, 	 -33, 	 -36, 	 -35, 	 -26, 	 -22, 		 -24, 	 -31, 	 -39, 	 -36, 	 -47, 	 -54, 	 -50, 	 -48, 	 -56, 	 -52, 	 -47, 	 -34, 	 -28, 	 -20, 	 -15, 	 -15, 	  11, 	  35, 	  24, 	  24, 	  41, 	  47, 	  62, 	  62, 	  66, 	  67, 	  59, 	  57, 	  59, 	  49, 	  54, 	  54, 	  48, 	  53, 	  57, 	  48, 	  53, 	  37, 	  20, 	  14, 	  15, 	  11, 	  38, 	  54, 	  48, 	  37, 	  10, 	 -56, 	 -61, 	 -49, 	 -46, 	 -47, 	 -58, 	 -60, 	 -63, 	 -68, 	 -68, 	 -73, 	 -76, 	 -77, 	 -77, 	 -82, 	 -79, 	 -81, 	
 -66, 	 -65, 	 -60, 	 -61, 	 -62, 	 -62, 	 -62, 	 -62, 	 -60, 	 -50, 	 -43, 	 -39, 	 -38, 	 -38, 	 -41, 	 -44, 	 -47, 	 -49, 	 -56, 	 -57, 	 -54, 	 -43, 	 -33, 	 -29, 	 -31, 	 -32, 	 -29, 	 -35, 	 -40, 	 -46, 	 -50, 	 -50, 	 -52, 	 -65, 	 -74, 	 -84, 	 -85, 	 -86, 	 -87, 	 -87, 	 -88, 	 -89, 	 -90, 	 -90, 	 -88, 	 -85, 	 -76, 	 -79, 	 -73, 	 -50, 	 -19, 	 -50, 	 -53, 	 -52, 	 -35, 	  16, 	  76, 	  -4, 	 -23, 	 -31, 	 -29, 	 -33, 	 -27, 	 -24, 		 -28, 	 -36, 	 -35, 	 -40, 	 -37, 	 -56, 	 -50, 	 -48, 	 -47, 	 -47, 	 -46, 	 -29, 	 -29, 	 -24, 	  -8, 	  20, 	   7, 	  28, 	  41, 	  31, 	  33, 	  38, 	  60, 	  62, 	  63, 	  65, 	  58, 	  51, 	  62, 	  52, 	  51, 	  55, 	  54, 	  52, 	  60, 	  48, 	  53, 	  53, 	  29, 	  17, 	  18, 	   5, 	  15, 	  55, 	  52, 	  45, 	  28, 	 -24, 	 -58, 	 -77, 	 -79, 	 -82, 	 -83, 	 -81, 	 -83, 	 -86, 	 -84, 	 -87, 	 -83, 	 -87, 	 -86, 	 -86, 	 -86, 	 -87, 	
 -68, 	 -65, 	 -60, 	 -62, 	 -63, 	 -62, 	 -64, 	 -64, 	 -66, 	 -61, 	 -52, 	 -45, 	 -43, 	 -43, 	 -44, 	 -45, 	 -45, 	 -42, 	 -45, 	 -51, 	 -59, 	 -53, 	 -44, 	 -37, 	 -35, 	 -36, 	 -32, 	 -35, 	 -39, 	 -47, 	 -51, 	 -50, 	 -52, 	 -58, 	 -74, 	 -82, 	 -86, 	 -85, 	 -86, 	 -86, 	 -86, 	 -89, 	 -88, 	 -89, 	 -90, 	 -88, 	 -76, 	 -80, 	 -79, 	 -73, 	 -36, 	 -36, 	 -53, 	 -52, 	 -35, 	   1, 	  80, 	  35, 	 -22, 	 -23, 	 -26, 	 -37, 	 -34, 	 -24, 		 -35, 	 -44, 	 -34, 	 -36, 	 -37, 	 -49, 	 -54, 	 -46, 	 -48, 	 -44, 	 -42, 	 -42, 	 -34, 	 -28, 	 -17, 	  43, 	  12, 	  20, 	  44, 	  44, 	  49, 	  43, 	  54, 	  63, 	  65, 	  63, 	  63, 	  47, 	  51, 	  63, 	  60, 	  50, 	  49, 	  52, 	  61, 	  55, 	  49, 	  52, 	  29, 	  28, 	  16, 	   5, 	   2, 	  36, 	  50, 	  46, 	  39, 	  -5, 	 -48, 	 -78, 	 -86, 	 -85, 	 -85, 	 -86, 	 -85, 	 -89, 	 -86, 	 -86, 	 -88, 	 -85, 	 -85, 	 -85, 	 -87, 	 -83, 	
 -69, 	 -69, 	 -67, 	 -64, 	 -65, 	 -64, 	 -62, 	 -61, 	 -67, 	 -66, 	 -64, 	 -55, 	 -50, 	 -44, 	 -43, 	 -46, 	 -48, 	 -46, 	 -43, 	 -45, 	 -48, 	 -58, 	 -49, 	 -42, 	 -40, 	 -41, 	 -37, 	 -35, 	 -38, 	 -46, 	 -51, 	 -51, 	 -50, 	 -51, 	 -67, 	 -82, 	 -88, 	 -84, 	 -85, 	 -86, 	 -85, 	 -88, 	 -87, 	 -88, 	 -90, 	 -90, 	 -83, 	 -80, 	 -77, 	 -77, 	 -58, 	 -29, 	 -48, 	 -47, 	   6, 	  23, 	  48, 	  82, 	 -16, 	 -26, 	 -26, 	 -26, 	 -32, 	 -31, 		 -37, 	 -40, 	 -31, 	 -33, 	 -32, 	 -39, 	 -52, 	 -49, 	 -48, 	 -52, 	 -46, 	 -44, 	 -36, 	 -26, 	 -18, 	  20, 	  15, 	  14, 	  36, 	  52, 	  54, 	  46, 	  53, 	  62, 	  63, 	  61, 	  66, 	  50, 	  42, 	  60, 	  57, 	  44, 	  46, 	  44, 	  57, 	  59, 	  43, 	  49, 	  34, 	  26, 	  18, 	   8, 	  -2, 	   4, 	  39, 	  46, 	  48, 	  34, 	   6, 	 -69, 	 -82, 	 -83, 	 -82, 	 -82, 	 -84, 	 -81, 	 -80, 	 -80, 	 -77, 	 -76, 	 -68, 	 -64, 	 -56, 	 -55, 	
 -68, 	 -67, 	 -68, 	 -67, 	 -65, 	 -65, 	 -66, 	 -62, 	 -65, 	 -66, 	 -69, 	 -63, 	 -59, 	 -54, 	 -48, 	 -47, 	 -48, 	 -49, 	 -44, 	 -41, 	 -42, 	 -49, 	 -56, 	 -48, 	 -43, 	 -44, 	 -40, 	 -39, 	 -39, 	 -41, 	 -47, 	 -54, 	 -50, 	 -48, 	 -52, 	 -73, 	 -84, 	 -84, 	 -83, 	 -86, 	 -86, 	 -84, 	 -88, 	 -91, 	 -89, 	 -89, 	 -90, 	 -80, 	 -79, 	 -78, 	 -73, 	 -41, 	 -32, 	 -36, 	  19, 	  11, 	  23, 	  96, 	   8, 	 -26, 	 -23, 	 -28, 	 -28, 	 -34, 		 -35, 	 -30, 	 -24, 	 -29, 	 -26, 	 -32, 	 -48, 	 -54, 	 -51, 	 -48, 	 -47, 	 -37, 	 -35, 	 -20, 	 -18, 	  -9, 	  10, 	   6, 	  32, 	  51, 	  49, 	  49, 	  57, 	  60, 	  61, 	  63, 	  63, 	  54, 	  37, 	  51, 	  61, 	  50, 	  47, 	  38, 	  47, 	  57, 	  46, 	  47, 	  40, 	  26, 	  24, 	  11, 	  -1, 	  -8, 	  25, 	  46, 	  49, 	  39, 	  29, 	 -21, 	 -21, 	 -37, 	 -44, 	 -34, 	 -36, 	 -36, 	 -21, 	 -14, 	 -12, 	  -6, 	   6, 	  29, 	   7, 	  -5, 	
 -71, 	 -70, 	 -69, 	 -71, 	 -69, 	 -66, 	 -67, 	 -65, 	 -68, 	 -69, 	 -69, 	 -68, 	 -64, 	 -60, 	 -58, 	 -57, 	 -55, 	 -53, 	 -51, 	 -41, 	 -40, 	 -42, 	 -51, 	 -52, 	 -49, 	 -44, 	 -39, 	 -40, 	 -40, 	 -44, 	 -45, 	 -49, 	 -50, 	 -46, 	 -44, 	 -53, 	 -79, 	 -80, 	 -84, 	 -85, 	 -84, 	 -84, 	 -87, 	 -85, 	 -88, 	 -91, 	 -89, 	 -83, 	 -77, 	 -79, 	 -77, 	 -60, 	 -23, 	 -36, 	 -21, 	 -26, 	  -9, 	  72, 	  48, 	 -26, 	 -32, 	 -29, 	 -35, 	 -32, 		 -35, 	 -39, 	 -29, 	 -20, 	 -22, 	 -29, 	 -38, 	 -48, 	 -45, 	 -25, 	 -41, 	 -43, 	 -31, 	 -20, 	 -15, 	 -16, 	   2, 	 -12, 	  23, 	  47, 	  55, 	  54, 	  52, 	  66, 	  59, 	  59, 	  62, 	  60, 	  51, 	  49, 	  61, 	  58, 	  48, 	  45, 	  40, 	  53, 	  49, 	  43, 	  45, 	  32, 	  23, 	  18, 	   4, 	   1, 	   7, 	  39, 	  45, 	  41, 	  17, 	  -6, 	  46, 	  46, 	  49, 	  36, 	  27, 	   5, 	 -28, 	 -33, 	 -45, 	 -43, 	 -44, 	 -19, 	 -20, 	 -32, 	
 -73, 	 -71, 	 -72, 	 -72, 	 -70, 	 -70, 	 -69, 	 -69, 	 -67, 	 -67, 	 -68, 	 -67, 	 -66, 	 -63, 	 -59, 	 -62, 	 -59, 	 -54, 	 -50, 	 -44, 	 -42, 	 -37, 	 -45, 	 -49, 	 -49, 	 -49, 	 -45, 	 -42, 	 -36, 	 -42, 	 -42, 	 -44, 	 -48, 	 -43, 	 -32, 	 -35, 	 -62, 	 -79, 	 -83, 	 -81, 	 -85, 	 -84, 	 -85, 	 -87, 	 -88, 	 -87, 	 -86, 	 -88, 	 -79, 	 -75, 	 -80, 	 -72, 	 -43, 	 -17, 	 -45, 	 -39, 	 -28, 	  33, 	  86, 	 -15, 	 -37, 	 -41, 	 -42, 	 -41, 		 -35, 	 -40, 	 -38, 	 -23, 	 -21, 	 -31, 	 -36, 	 -41, 	 -42, 	 -21, 	 -31, 	 -25, 	 -28, 	 -14, 	 -14, 	 -16, 	 -10, 	  -9, 	   3, 	  33, 	  47, 	  48, 	  57, 	  66, 	  60, 	  53, 	  53, 	  55, 	  50, 	  37, 	  47, 	  53, 	  50, 	  51, 	  43, 	  55, 	  59, 	  47, 	  48, 	  42, 	  27, 	  22, 	  16, 	  19, 	   4, 	  29, 	  44, 	  45, 	  33, 	  -6, 	  41, 	  46, 	  47, 	  50, 	  40, 	  16, 	 -37, 	 -42, 	 -20, 	 -48, 	 -50, 	 -53, 	 -40, 	 -35, 	
 -77, 	 -75, 	 -76, 	 -73, 	 -72, 	 -72, 	 -71, 	 -68, 	 -69, 	 -68, 	 -69, 	 -68, 	 -67, 	 -64, 	 -61, 	 -61, 	 -63, 	 -57, 	 -53, 	 -46, 	 -41, 	 -36, 	 -37, 	 -42, 	 -49, 	 -52, 	 -49, 	 -45, 	 -38, 	 -37, 	 -38, 	 -40, 	 -40, 	 -38, 	 -30, 	 -30, 	 -37, 	 -68, 	 -80, 	 -82, 	 -83, 	 -84, 	 -83, 	 -87, 	 -85, 	 -87, 	 -88, 	 -89, 	 -83, 	 -73, 	 -76, 	 -76, 	 -62, 	 -18, 	 -32, 	 -38, 	 -34, 	   1, 	  90, 	  32, 	 -32, 	 -42, 	 -42, 	 -38, 		 -37, 	 -37, 	 -40, 	 -32, 	 -36, 	 -32, 	 -30, 	 -41, 	 -40, 	 -24, 	 -13, 	  -1, 	  -9, 	 -18, 	  -7, 	   3, 	  -1, 	   1, 	 -13, 	  28, 	  31, 	  32, 	  48, 	  63, 	  60, 	  58, 	  46, 	  44, 	  52, 	  45, 	  45, 	  51, 	  48, 	  39, 	  45, 	  54, 	  58, 	  46, 	  51, 	  49, 	  38, 	  29, 	  24, 	  12, 	  17, 	  17, 	  45, 	  50, 	  38, 	  -3, 	 -28, 	  17, 	  28, 	  28, 	 -20, 	 -40, 	 -40, 	 -51, 	 -49, 	 -41, 	 -56, 	 -50, 	 -39, 	 -13, 	
 -80, 	 -80, 	 -79, 	 -75, 	 -78, 	 -72, 	 -73, 	 -71, 	 -70, 	 -70, 	 -68, 	 -67, 	 -67, 	 -66, 	 -63, 	 -61, 	 -62, 	 -57, 	 -49, 	 -47, 	 -41, 	 -33, 	 -33, 	 -36, 	 -41, 	 -51, 	 -56, 	 -49, 	 -45, 	 -34, 	 -33, 	 -35, 	 -37, 	 -34, 	 -32, 	 -21, 	 -26, 	 -48, 	 -76, 	 -81, 	 -82, 	 -84, 	 -84, 	 -84, 	 -82, 	 -86, 	 -88, 	 -88, 	 -88, 	 -73, 	 -73, 	 -76, 	 -75, 	 -42, 	 -12, 	 -40, 	 -34, 	 -13, 	  64, 	  85, 	 -26, 	 -36, 	 -29, 	 -16, 		 -24, 	 -29, 	 -35, 	 -36, 	 -32, 	 -29, 	 -32, 	 -42, 	 -37, 	 -24, 	   2, 	  14, 	   9, 	  -4, 	 -13, 	  11, 	  20, 	  21, 	   3, 	   1, 	  36, 	  34, 	  50, 	  56, 	  55, 	  60, 	  48, 	  55, 	  53, 	  48, 	  42, 	  43, 	  41, 	  27, 	  40, 	  52, 	  46, 	  45, 	  48, 	  48, 	  42, 	  37, 	  23, 	  15, 	  25, 	   2, 	  24, 	  47, 	  40, 	  28, 	 -10, 	   6, 	   6, 	   9, 	 -35, 	 -61, 	 -43, 	 -48, 	 -62, 	 -44, 	 -51, 	 -51, 	 -33, 	 -22, 	
 -82, 	 -81, 	 -79, 	 -80, 	 -78, 	 -78, 	 -73, 	 -73, 	 -74, 	 -72, 	 -70, 	 -69, 	 -68, 	 -69, 	 -66, 	 -64, 	 -62, 	 -60, 	 -52, 	 -44, 	 -42, 	 -31, 	 -35, 	 -33, 	 -37, 	 -45, 	 -55, 	 -57, 	 -48, 	 -41, 	 -27, 	 -33, 	 -27, 	 -27, 	 -27, 	 -21, 	 -21, 	 -29, 	 -59, 	 -78, 	 -81, 	 -83, 	 -82, 	 -81, 	 -82, 	 -88, 	 -84, 	 -89, 	 -89, 	 -82, 	 -77, 	 -75, 	 -76, 	 -63, 	 -16, 	 -18, 	 -21, 	 -18, 	  45, 	  99, 	  21, 	 -35, 	 -23, 	 -14, 		 -20, 	 -21, 	 -32, 	 -29, 	   2, 	 -21, 	 -29, 	 -31, 	 -33, 	 -18, 	 -24, 	  11, 	  23, 	  -2, 	  11, 	  16, 	  21, 	  56, 	  27, 	 -13, 	   7, 	  36, 	  46, 	  49, 	  50, 	  57, 	  46, 	  53, 	  55, 	  53, 	  49, 	  47, 	  48, 	  36, 	  31, 	  45, 	  39, 	  51, 	  44, 	  53, 	  43, 	  31, 	  33, 	  21, 	   9, 	  -7, 	   0, 	  31, 	  38, 	  34, 	  11, 	  17, 	   2, 	 -48, 	 -61, 	 -78, 	 -63, 	 -37, 	 -30, 	 -43, 	 -46, 	 -34, 	 -22, 	 -15, 	
 -83, 	 -85, 	 -85, 	 -80, 	 -80, 	 -79, 	 -77, 	 -75, 	 -73, 	 -70, 	 -72, 	 -72, 	 -69, 	 -69, 	 -65, 	 -66, 	 -63, 	 -60, 	 -55, 	 -46, 	 -36, 	 -31, 	 -33, 	 -33, 	 -33, 	 -41, 	 -47, 	 -59, 	 -60, 	 -48, 	 -36, 	 -25, 	 -26, 	 -24, 	 -20, 	 -21, 	 -20, 	 -23, 	 -36, 	 -68, 	 -78, 	 -77, 	 -79, 	 -78, 	 -82, 	 -85, 	 -84, 	 -87, 	 -87, 	 -88, 	 -76, 	 -68, 	 -75, 	 -69, 	 -44, 	  -9, 	 -18, 	 -17, 	  16, 	  90, 	  71, 	 -22, 	 -36, 	 -14, 		 -16, 	 -14, 	 -30, 	  -6, 	  12, 	 -12, 	 -18, 	 -17, 	 -27, 	 -26, 	 -24, 	  13, 	  41, 	  24, 	  13, 	  26, 	  45, 	  35, 	  38, 	   8, 	  -9, 	  35, 	  40, 	  26, 	  32, 	  25, 	  11, 	  30, 	  47, 	  44, 	  50, 	  51, 	  47, 	  41, 	  34, 	  39, 	  44, 	  47, 	  49, 	  47, 	  49, 	  32, 	  29, 	  37, 	   4, 	   4, 	  -2, 	  20, 	  43, 	  43, 	  22, 	   8, 	   5, 	  -6, 	 -41, 	 -70, 	 -50, 	  -5, 	  22, 	  26, 	  -8, 	 -23, 	 -18, 	  -1, 	
 -84, 	 -84, 	 -85, 	 -85, 	 -85, 	 -81, 	 -79, 	 -79, 	 -78, 	 -76, 	 -72, 	 -73, 	 -70, 	 -67, 	 -66, 	 -65, 	 -65, 	 -62, 	 -59, 	 -52, 	 -38, 	 -32, 	 -31, 	 -33, 	 -37, 	 -39, 	 -42, 	 -53, 	 -65, 	 -54, 	 -44, 	 -28, 	 -23, 	 -22, 	 -22, 	 -20, 	 -17, 	 -21, 	 -26, 	 -45, 	 -68, 	 -73, 	 -71, 	 -73, 	 -77, 	 -82, 	 -88, 	 -88, 	 -86, 	 -87, 	 -83, 	 -64, 	 -73, 	 -73, 	 -62, 	 -21, 	  -5, 	 -21, 	 -10, 	  66, 	  99, 	  -5, 	 -34, 	 -19, 		 -18, 	 -10, 	 -18, 	   0, 	   6, 	  -7, 	 -10, 	 -18, 	 -14, 	 -27, 	   8, 	   5, 	  47, 	  30, 	  34, 	  15, 	  29, 	  34, 	  49, 	  28, 	  15, 	  31, 	  42, 	  17, 	  -4, 	  12, 	  16, 	  23, 	  11, 	  42, 	  52, 	  45, 	  51, 	  43, 	  36, 	  36, 	  52, 	  53, 	  55, 	  46, 	  50, 	  33, 	  27, 	  37, 	  24, 	  13, 	  20, 	  14, 	  47, 	  44, 	  33, 	   4, 	  17, 	  -2, 	 -21, 	 -35, 	 -31, 	 -26, 	 -26, 	   8, 	  21, 	  37, 	  18, 	  22, 	
 -84, 	 -84, 	 -84, 	 -85, 	 -83, 	 -83, 	 -84, 	 -81, 	 -79, 	 -77, 	 -73, 	 -73, 	 -72, 	 -71, 	 -68, 	 -65, 	 -63, 	 -66, 	 -62, 	 -57, 	 -49, 	 -34, 	 -31, 	 -35, 	 -38, 	 -42, 	 -38, 	 -48, 	 -59, 	 -63, 	 -47, 	 -36, 	 -21, 	 -20, 	 -20, 	 -18, 	 -19, 	 -19, 	 -27, 	 -30, 	 -54, 	 -67, 	 -66, 	 -65, 	 -71, 	 -84, 	 -84, 	 -84, 	 -88, 	 -90, 	 -89, 	 -72, 	 -71, 	 -74, 	 -69, 	 -47, 	   4, 	 -22, 	 -16, 	  40, 	  98, 	  31, 	 -37, 	 -35, 		 -26, 	 -24, 	 -18, 	  -3, 	  -8, 	 -10, 	 -13, 	  -8, 	 -12, 	 -16, 	  -5, 	  14, 	  20, 	  28, 	  31, 	  17, 	  34, 	  33, 	  29, 	  41, 	  24, 	  21, 	  40, 	  14, 	   1, 	  14, 	  52, 	  52, 	  15, 	  31, 	  51, 	  42, 	  42, 	  45, 	  39, 	  41, 	  49, 	  53, 	  55, 	  52, 	  50, 	  36, 	  31, 	  34, 	  30, 	  18, 	  56, 	  18, 	  39, 	  42, 	  41, 	  11, 	 -12, 	 -28, 	 -39, 	 -20, 	 -44, 	 -45, 	 -53, 	 -52, 	 -45, 	 -18, 	   7, 	  21, 	
 -87, 	 -85, 	 -85, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -83, 	 -81, 	 -77, 	 -75, 	 -73, 	 -72, 	 -69, 	 -68, 	 -66, 	 -62, 	 -64, 	 -60, 	 -58, 	 -49, 	 -35, 	 -37, 	 -41, 	 -41, 	 -42, 	 -49, 	 -57, 	 -59, 	 -56, 	 -42, 	 -30, 	 -17, 	 -20, 	 -21, 	 -18, 	 -16, 	 -25, 	 -29, 	 -37, 	 -59, 	 -63, 	 -59, 	 -60, 	 -71, 	 -83, 	 -88, 	 -87, 	 -91, 	 -90, 	 -85, 	 -74, 	 -76, 	 -76, 	 -65, 	 -10, 	  -8, 	 -17, 	  22, 	  90, 	  76, 	 -29, 	 -42, 		 -39, 	 -37, 	 -14, 	 -11, 	 -17, 	 -20, 	 -18, 	  -4, 	  -8, 	 -14, 	 -17, 	  23, 	   1, 	  43, 	  15, 	  12, 	  28, 	  37, 	  44, 	  55, 	  32, 	  21, 	  38, 	  34, 	  11, 	  45, 	  53, 	  59, 	  37, 	  26, 	  44, 	  33, 	  29, 	  43, 	  40, 	  35, 	  43, 	  47, 	  55, 	  49, 	  50, 	  51, 	  32, 	  31, 	  41, 	  26, 	  43, 	  39, 	  28, 	  42, 	  33, 	  25, 	 -21, 	 -53, 	 -53, 	 -37, 	 -61, 	 -62, 	 -78, 	 -79, 	 -49, 	 -43, 	 -45, 	 -50, 	
 -89, 	 -88, 	 -87, 	 -86, 	 -85, 	 -84, 	 -84, 	 -84, 	 -84, 	 -83, 	 -79, 	 -75, 	 -73, 	 -72, 	 -69, 	 -71, 	 -68, 	 -66, 	 -65, 	 -65, 	 -63, 	 -56, 	 -50, 	 -41, 	 -45, 	 -47, 	 -46, 	 -47, 	 -51, 	 -56, 	 -60, 	 -52, 	 -39, 	 -27, 	 -19, 	 -24, 	 -17, 	 -19, 	 -25, 	 -34, 	 -32, 	 -52, 	 -60, 	 -60, 	 -56, 	 -57, 	 -82, 	 -88, 	 -89, 	 -91, 	 -90, 	 -90, 	 -83, 	 -78, 	 -76, 	 -73, 	 -42, 	   5, 	 -17, 	  13, 	  72, 	  97, 	  15, 	 -39, 		 -42, 	 -34, 	 -26, 	 -24, 	 -28, 	 -27, 	  -9, 	  -3, 	  -6, 	  -9, 	 -26, 	   0, 	  11, 	  22, 	  43, 	  12, 	   9, 	   8, 	  26, 	  46, 	  22, 	  23, 	  28, 	  49, 	  44, 	  54, 	  50, 	  55, 	  30, 	   8, 	  27, 	  19, 	   9, 	  43, 	  36, 	  28, 	  31, 	  39, 	  53, 	  46, 	  37, 	  47, 	  50, 	  42, 	  32, 	  38, 	  33, 	  42, 	  21, 	  29, 	  37, 	  25, 	 -37, 	 -59, 	 -48, 	 -42, 	 -58, 	 -79, 	 -70, 	 -72, 	 -44, 	 -50, 	 -59, 	 -52, 	
 -83, 	 -86, 	 -88, 	 -89, 	 -85, 	 -84, 	 -84, 	 -84, 	 -83, 	 -83, 	 -83, 	 -81, 	 -77, 	 -75, 	 -72, 	 -70, 	 -70, 	 -68, 	 -67, 	 -64, 	 -64, 	 -61, 	 -62, 	 -51, 	 -48, 	 -49, 	 -50, 	 -47, 	 -49, 	 -52, 	 -55, 	 -53, 	 -47, 	 -32, 	 -22, 	 -20, 	 -24, 	 -19, 	 -23, 	 -32, 	 -37, 	 -42, 	 -56, 	 -56, 	 -51, 	 -52, 	 -72, 	 -87, 	 -89, 	 -91, 	 -89, 	 -91, 	 -88, 	 -79, 	 -75, 	 -73, 	 -61, 	 -15, 	  -7, 	   7, 	  51, 	  95, 	  62, 	 -35, 		 -34, 	 -27, 	 -26, 	 -28, 	 -23, 	 -14, 	   3, 	   1, 	  -3, 	 -15, 	 -26, 	  -6, 	  12, 	   7, 	  23, 	   7, 	   3, 	  14, 	  32, 	  43, 	  18, 	  17, 	  17, 	  48, 	  49, 	  50, 	  52, 	  53, 	  26, 	  13, 	   3, 	  -3, 	   3, 	  44, 	  45, 	  43, 	  38, 	  38, 	  43, 	  43, 	  28, 	  28, 	  38, 	  44, 	  37, 	  33, 	  32, 	  25, 	  20, 	  15, 	  34, 	  24, 	   4, 	 -42, 	 -37, 	 -37, 	 -46, 	 -76, 	 -82, 	 -74, 	 -44, 	 -44, 	 -36, 	 -71, 	
 -85, 	 -82, 	 -84, 	 -86, 	 -90, 	 -88, 	 -86, 	 -85, 	 -86, 	 -83, 	 -84, 	 -83, 	 -81, 	 -79, 	 -74, 	 -71, 	 -70, 	 -69, 	 -70, 	 -68, 	 -62, 	 -65, 	 -67, 	 -62, 	 -55, 	 -51, 	 -53, 	 -51, 	 -47, 	 -50, 	 -50, 	 -55, 	 -53, 	 -39, 	 -29, 	 -24, 	 -24, 	 -25, 	 -24, 	 -30, 	 -37, 	 -39, 	 -48, 	 -52, 	 -49, 	 -49, 	 -59, 	 -85, 	 -88, 	 -89, 	 -91, 	 -91, 	 -91, 	 -84, 	 -81, 	 -74, 	 -69, 	 -50, 	   0, 	   8, 	  36, 	  89, 	  91, 	 -14, 		 -34, 	 -27, 	 -21, 	 -21, 	 -10, 	  -3, 	   7, 	  10, 	  -2, 	 -16, 	 -21, 	 -27, 	  16, 	  10, 	  17, 	   9, 	  -9, 	  10, 	  46, 	  23, 	  -2, 	  12, 	   1, 	  21, 	  48, 	  50, 	  53, 	  54, 	  36, 	  22, 	  14, 	 -20, 	  -8, 	  37, 	  44, 	  42, 	  39, 	  41, 	  30, 	  13, 	  23, 	  10, 	  26, 	  33, 	  45, 	  34, 	  31, 	  19, 	   3, 	  -5, 	  15, 	  25, 	  23, 	 -33, 	 -33, 	 -40, 	 -55, 	 -65, 	 -60, 	 -70, 	 -43, 	 -27, 	 -44, 	 -67, 	
 -81, 	 -83, 	 -82, 	 -83, 	 -83, 	 -86, 	 -89, 	 -87, 	 -85, 	 -83, 	 -84, 	 -83, 	 -83, 	 -81, 	 -77, 	 -74, 	 -72, 	 -73, 	 -70, 	 -68, 	 -68, 	 -66, 	 -69, 	 -64, 	 -63, 	 -56, 	 -49, 	 -52, 	 -49, 	 -48, 	 -50, 	 -49, 	 -50, 	 -47, 	 -40, 	 -29, 	 -31, 	 -25, 	 -23, 	 -29, 	 -34, 	 -42, 	 -48, 	 -53, 	 -49, 	 -52, 	 -56, 	 -75, 	 -87, 	 -89, 	 -89, 	 -91, 	 -90, 	 -86, 	 -80, 	 -75, 	 -75, 	 -65, 	 -24, 	  12, 	  29, 	  66, 	  94, 	  17, 		 -40, 	 -26, 	 -27, 	 -22, 	  -8, 	   0, 	   4, 	  -1, 	   3, 	  -6, 	 -21, 	 -26, 	   4, 	  13, 	   9, 	  20, 	   2, 	 -13, 	  33, 	  15, 	   3, 	   6, 	  10, 	  19, 	  38, 	  43, 	  47, 	  45, 	  28, 	  28, 	  25, 	 -14, 	 -17, 	  12, 	  36, 	  34, 	  30, 	  23, 	  21, 	  23, 	  17, 	   4, 	   2, 	  19, 	  40, 	  14, 	  10, 	  19, 	   4, 	 -25, 	 -12, 	  16, 	  30, 	 -24, 	 -44, 	 -49, 	 -40, 	 -28, 	 -52, 	 -49, 	 -45, 	 -20, 	 -56, 	 -74, 	
 -81, 	 -82, 	 -81, 	 -82, 	 -83, 	 -84, 	 -85, 	 -87, 	 -87, 	 -86, 	 -85, 	 -85, 	 -83, 	 -85, 	 -82, 	 -79, 	 -75, 	 -72, 	 -70, 	 -72, 	 -70, 	 -66, 	 -67, 	 -66, 	 -65, 	 -59, 	 -56, 	 -48, 	 -49, 	 -50, 	 -46, 	 -49, 	 -47, 	 -50, 	 -44, 	 -37, 	 -31, 	 -28, 	 -27, 	 -27, 	 -34, 	 -42, 	 -48, 	 -58, 	 -61, 	 -56, 	 -63, 	 -70, 	 -85, 	 -88, 	 -89, 	 -89, 	 -90, 	 -89, 	 -81, 	 -72, 	 -77, 	 -71, 	 -43, 	   7, 	  27, 	  62, 	  92, 	  38, 		 -31, 	 -34, 	 -21, 	 -17, 	  -6, 	  -5, 	   7, 	  -8, 	   7, 	   1, 	 -20, 	  -7, 	 -14, 	  -8, 	  -9, 	   2, 	  -5, 	 -20, 	   1, 	  12, 	  -6, 	 -11, 	   4, 	  20, 	  27, 	  35, 	  44, 	  46, 	  13, 	   6, 	  11, 	 -20, 	 -21, 	  -5, 	  25, 	  23, 	  25, 	  24, 	  24, 	  28, 	   2, 	 -15, 	 -30, 	 -20, 	   7, 	 -10, 	 -29, 	 -13, 	  -6, 	 -37, 	 -34, 	  12, 	  25, 	  -2, 	 -55, 	 -61, 	 -43, 	 -12, 	 -16, 	   6, 	 -24, 	 -16, 	 -48, 	 -75, 	
 -82, 	 -82, 	 -81, 	 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -85, 	 -85, 	 -86, 	 -84, 	 -84, 	 -84, 	 -83, 	 -83, 	 -77, 	 -74, 	 -70, 	 -72, 	 -71, 	 -68, 	 -68, 	 -67, 	 -66, 	 -63, 	 -55, 	 -50, 	 -47, 	 -50, 	 -49, 	 -43, 	 -48, 	 -46, 	 -51, 	 -42, 	 -34, 	 -32, 	 -29, 	 -31, 	 -35, 	 -45, 	 -54, 	 -59, 	 -65, 	 -66, 	 -63, 	 -68, 	 -80, 	 -88, 	 -89, 	 -90, 	 -87, 	 -91, 	 -89, 	 -81, 	 -76, 	 -75, 	 -62, 	 -13, 	  21, 	  58, 	  94, 	  76, 		 -23, 	 -36, 	 -26, 	 -25, 	 -25, 	 -16, 	 -17, 	   2, 	   8, 	   6, 	  -9, 	  -6, 	 -18, 	 -23, 	 -17, 	 -18, 	 -16, 	 -23, 	 -21, 	   1, 	 -41, 	 -20, 	 -11, 	  11, 	  22, 	  39, 	  40, 	  19, 	  21, 	   7, 	   0, 	 -15, 	 -12, 	  -9, 	  30, 	  29, 	  22, 	  25, 	  24, 	  22, 	 -10, 	 -24, 	 -38, 	 -41, 	 -24, 	 -15, 	 -28, 	 -29, 	 -26, 	 -39, 	 -35, 	 -11, 	  23, 	  19, 	 -44, 	 -58, 	 -41, 	 -25, 	 -14, 	 -11, 	  30, 	  21, 	 -23, 	 -58, 	
 -85, 	 -85, 	 -85, 	 -84, 	 -85, 	 -84, 	 -84, 	 -82, 	 -83, 	 -83, 	 -87, 	 -88, 	 -83, 	 -85, 	 -84, 	 -86, 	 -81, 	 -79, 	 -76, 	 -74, 	 -73, 	 -69, 	 -70, 	 -68, 	 -68, 	 -67, 	 -60, 	 -54, 	 -51, 	 -47, 	 -48, 	 -45, 	 -42, 	 -46, 	 -49, 	 -47, 	 -43, 	 -35, 	 -35, 	 -31, 	 -39, 	 -47, 	 -52, 	 -62, 	 -65, 	 -70, 	 -70, 	 -73, 	 -78, 	 -87, 	 -88, 	 -91, 	 -88, 	 -89, 	 -90, 	 -91, 	 -88, 	 -83, 	 -73, 	 -38, 	   6, 	  37, 	  91, 	  89, 		  -5, 	 -33, 	 -38, 	 -37, 	 -36, 	 -34, 	 -32, 	  -9, 	  -9, 	  -1, 	 -14, 	 -17, 	  -5, 	 -20, 	 -29, 	 -21, 	 -22, 	 -27, 	 -35, 	 -14, 	 -47, 	 -31, 	 -22, 	   6, 	  26, 	  38, 	  17, 	   0, 	   1, 	  -3, 	 -15, 	 -27, 	 -10, 	 -22, 	  -5, 	 -11, 	 -18, 	  -3, 	 -28, 	 -24, 	 -33, 	 -54, 	 -61, 	 -61, 	 -57, 	 -49, 	 -63, 	 -65, 	 -67, 	 -68, 	 -67, 	 -57, 	 -28, 	  -4, 	 -28, 	 -66, 	 -56, 	 -54, 	 -39, 	 -31, 	  -7, 	  16, 	  34, 	  35, 	
 -86, 	 -86, 	 -87, 	 -87, 	 -86, 	 -87, 	 -86, 	 -84, 	 -83, 	 -83, 	 -85, 	 -86, 	 -87, 	 -84, 	 -83, 	 -84, 	 -84, 	 -84, 	 -79, 	 -75, 	 -73, 	 -70, 	 -72, 	 -68, 	 -67, 	 -69, 	 -66, 	 -57, 	 -54, 	 -46, 	 -48, 	 -46, 	 -41, 	 -43, 	 -47, 	 -52, 	 -46, 	 -42, 	 -39, 	 -37, 	 -39, 	 -45, 	 -54, 	 -68, 	 -68, 	 -70, 	 -73, 	 -77, 	 -81, 	 -85, 	 -89, 	 -89, 	 -88, 	 -89, 	 -91, 	 -89, 	 -91, 	 -87, 	 -83, 	 -63, 	  -9, 	  20, 	  42, 	  59, 		 -29, 	 -50, 	 -44, 	 -46, 	 -45, 	 -50, 	 -48, 	 -39, 	 -37, 	 -38, 	 -41, 	 -39, 	 -27, 	 -42, 	 -60, 	 -50, 	 -38, 	 -49, 	 -54, 	 -58, 	 -71, 	 -57, 	 -54, 	 -52, 	 -45, 	 -55, 	 -63, 	 -65, 	 -67, 	 -72, 	 -71, 	 -75, 	 -74, 	 -75, 	 -76, 	 -81, 	 -78, 	 -79, 	 -82, 	 -78, 	 -77, 	 -82, 	 -80, 	 -83, 	 -81, 	 -81, 	 -83, 	 -79, 	 -78, 	 -83, 	 -86, 	 -83, 	 -80, 	 -73, 	 -54, 	 -68, 	 -63, 	 -64, 	 -69, 	 -65, 	 -48, 	 -40, 	 -36, 	 -19, 	
 -86, 	 -86, 	 -86, 	 -87, 	 -87, 	 -87, 	 -87, 	 -87, 	 -85, 	 -84, 	 -84, 	 -82, 	 -86, 	 -85, 	 -84, 	 -84, 	 -82, 	 -83, 	 -81, 	 -79, 	 -76, 	 -72, 	 -71, 	 -68, 	 -66, 	 -65, 	 -65, 	 -60, 	 -52, 	 -51, 	 -49, 	 -48, 	 -39, 	 -41, 	 -42, 	 -50, 	 -51, 	 -43, 	 -44, 	 -37, 	 -35, 	 -47, 	 -60, 	 -66, 	 -69, 	 -66, 	 -73, 	 -79, 	 -83, 	 -87, 	 -86, 	 -90, 	 -88, 	 -88, 	 -90, 	 -89, 	 -92, 	 -90, 	 -89, 	 -86, 	 -77, 	 -66, 	 -73, 	 -76, 		 -77, 	 -80, 	 -77, 	 -75, 	 -75, 	 -70, 	 -76, 	 -78, 	 -81, 	 -76, 	 -77, 	 -74, 	 -69, 	 -79, 	 -81, 	 -80, 	 -71, 	 -74, 	 -81, 	 -80, 	 -82, 	 -78, 	 -77, 	 -75, 	 -78, 	 -83, 	 -85, 	 -84, 	 -86, 	 -87, 	 -85, 	 -87, 	 -87, 	 -89, 	 -90, 	 -90, 	 -90, 	 -89, 	 -89, 	 -89, 	 -86, 	 -76, 	 -65, 	 -55, 	 -38, 	 -42, 	 -42, 	 -54, 	 -80, 	 -83, 	 -82, 	 -83, 	 -82, 	 -78, 	 -73, 	 -70, 	 -79, 	 -62, 	 -68, 	 -10, 	 -18, 	 -64, 	 -80, 	 -81, 	
 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -85, 	 -87, 	 -85, 	 -86, 	 -84, 	 -83, 	 -84, 	 -84, 	 -85, 	 -84, 	 -85, 	 -84, 	 -81, 	 -76, 	 -74, 	 -73, 	 -70, 	 -69, 	 -65, 	 -64, 	 -63, 	 -56, 	 -54, 	 -51, 	 -47, 	 -45, 	 -40, 	 -40, 	 -48, 	 -53, 	 -45, 	 -42, 	 -39, 	 -39, 	 -53, 	 -60, 	 -65, 	 -66, 	 -63, 	 -66, 	 -83, 	 -85, 	 -85, 	 -86, 	 -87, 	 -87, 	 -87, 	 -88, 	 -88, 	 -89, 	 -89, 	 -89, 	 -87, 	 -89, 	 -89, 	 -89, 	 -86, 		 -89, 	 -91, 	 -90, 	 -89, 	 -88, 	 -88, 	 -90, 	 -88, 	 -88, 	 -90, 	 -90, 	 -91, 	 -87, 	 -90, 	 -88, 	 -90, 	 -83, 	 -87, 	 -89, 	 -90, 	 -91, 	 -91, 	 -88, 	 -91, 	 -91, 	 -88, 	 -93, 	 -91, 	 -90, 	 -89, 	 -89, 	 -90, 	 -91, 	 -91, 	 -90, 	 -90, 	 -91, 	 -90, 	 -91, 	 -89, 	 -87, 	 -82, 	 -67, 	 -54, 	 -27, 	 -17, 	 -15, 	 -15, 	 -71, 	 -73, 	 -71, 	 -80, 	 -78, 	 -71, 	 -50, 	 -63, 	 -83, 	 -63, 	 -51, 	   2, 	  10, 	 -50, 	 -54, 	 -81, 	
 -85, 	 -85, 	 -85, 	 -85, 	 -85, 	 -85, 	 -86, 	 -86, 	 -85, 	 -86, 	 -86, 	 -86, 	 -81, 	 -84, 	 -84, 	 -87, 	 -86, 	 -85, 	 -84, 	 -83, 	 -81, 	 -78, 	 -74, 	 -71, 	 -68, 	 -68, 	 -67, 	 -68, 	 -60, 	 -57, 	 -54, 	 -48, 	 -44, 	 -40, 	 -36, 	 -47, 	 -52, 	 -49, 	 -45, 	 -41, 	 -44, 	 -49, 	 -57, 	 -63, 	 -62, 	 -59, 	 -57, 	 -74, 	 -83, 	 -83, 	 -83, 	 -86, 	 -88, 	 -86, 	 -89, 	 -87, 	 -89, 	 -90, 	 -90, 	 -91, 	 -89, 	 -89, 	 -89, 	 -90, 		 -91, 	 -89, 	 -90, 	 -93, 	 -92, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -89, 	 -92, 	 -91, 	 -91, 	 -91, 	 -92, 	 -84, 	 -90, 	 -91, 	 -92, 	 -91, 	 -91, 	 -91, 	 -92, 	 -91, 	 -91, 	 -90, 	 -93, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -90, 	 -90, 	 -92, 	 -85, 	 -67, 	 -54, 	 -32, 	 -11, 	 -16, 	  -6, 	 -64, 	 -76, 	 -74, 	 -79, 	 -78, 	 -62, 	 -55, 	 -60, 	 -77, 	 -65, 	 -33, 	 -54, 	 -29, 	 -48, 	   7, 	 -11, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -86, 	 -84, 	 -85, 	 -85, 	 -87, 	 -86, 	 -83, 	 -81, 	 -83, 	 -87, 	 -86, 	 -84, 	 -85, 	 -83, 	 -78, 	 -76, 	 -74, 	 -71, 	 -65, 	 -69, 	 -67, 	 -61, 	 -57, 	 -54, 	 -52, 	 -45, 	 -42, 	 -36, 	 -38, 	 -49, 	 -53, 	 -44, 	 -40, 	 -42, 	 -48, 	 -56, 	 -57, 	 -60, 	 -59, 	 -52, 	 -62, 	 -82, 	 -81, 	 -85, 	 -84, 	 -85, 	 -87, 	 -86, 	 -87, 	 -88, 	 -88, 	 -90, 	 -91, 	 -89, 	 -90, 	 -90, 	 -90, 		 -90, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -91, 	 -92, 	 -90, 	 -92, 	 -91, 	 -89, 	 -92, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -91, 	 -91, 	 -92, 	 -92, 	 -91, 	 -92, 	 -92, 	 -93, 	 -92, 	 -92, 	 -92, 	 -93, 	 -87, 	 -69, 	 -52, 	 -41, 	 -16, 	 -13, 	 -11, 	 -49, 	 -78, 	 -76, 	 -77, 	 -75, 	 -77, 	 -71, 	 -67, 	 -74, 	 -64, 	 -29, 	 -57, 	 -56, 	 -69, 	 -10, 	  35, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -85, 	 -85, 	 -85, 	 -84, 	 -85, 	 -85, 	 -84, 	 -82, 	 -82, 	 -85, 	 -88, 	 -84, 	 -83, 	 -85, 	 -81, 	 -77, 	 -74, 	 -71, 	 -66, 	 -68, 	 -65, 	 -62, 	 -57, 	 -54, 	 -53, 	 -46, 	 -38, 	 -38, 	 -39, 	 -44, 	 -51, 	 -51, 	 -43, 	 -40, 	 -43, 	 -49, 	 -54, 	 -54, 	 -54, 	 -45, 	 -45, 	 -73, 	 -80, 	 -82, 	 -85, 	 -84, 	 -85, 	 -86, 	 -86, 	 -88, 	 -88, 	 -89, 	 -91, 	 -90, 	 -90, 	 -90, 	 -89, 		 -90, 	 -90, 	 -90, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -91, 	 -91, 	 -91, 	 -91, 	 -90, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -91, 	 -91, 	 -91, 	 -92, 	 -90, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -92, 	 -92, 	 -87, 	 -77, 	 -64, 	 -46, 	 -17, 	  -9, 	 -13, 	 -36, 	 -81, 	 -85, 	 -84, 	 -86, 	 -89, 	 -84, 	 -75, 	 -82, 	 -67, 	 -28, 	 -66, 	 -64, 	 -72, 	 -47, 	   2, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -82, 	 -85, 	 -85, 	 -85, 	 -85, 	 -84, 	 -85, 	 -83, 	 -83, 	 -82, 	 -84, 	 -85, 	 -82, 	 -85, 	 -82, 	 -81, 	 -74, 	 -72, 	 -68, 	 -67, 	 -63, 	 -59, 	 -61, 	 -56, 	 -52, 	 -48, 	 -45, 	 -40, 	 -37, 	 -37, 	 -45, 	 -54, 	 -48, 	 -38, 	 -37, 	 -43, 	 -47, 	 -48, 	 -50, 	 -40, 	 -34, 	 -55, 	 -78, 	 -80, 	 -82, 	 -81, 	 -84, 	 -85, 	 -86, 	 -88, 	 -87, 	 -88, 	 -90, 	 -89, 	 -89, 	 -90, 	 -89, 		 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -91, 	 -91, 	 -92, 	 -91, 	 -92, 	 -91, 	 -92, 	 -90, 	 -92, 	 -92, 	 -91, 	 -91, 	 -90, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -91, 	 -90, 	 -90, 	 -91, 	 -91, 	 -90, 	 -92, 	 -92, 	 -92, 	 -92, 	 -93, 	 -93, 	 -91, 	 -90, 	 -82, 	 -67, 	 -49, 	 -28, 	 -10, 	 -15, 	 -25, 	 -79, 	 -80, 	 -81, 	 -81, 	 -84, 	 -87, 	 -90, 	 -86, 	 -75, 	 -33, 	 -60, 	 -54, 	 -56, 	 -67, 	 -33, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -85, 	 -85, 	 -83, 	 -85, 	 -87, 	 -85, 	 -84, 	 -85, 	 -84, 	 -85, 	 -81, 	 -83, 	 -87, 	 -84, 	 -83, 	 -83, 	 -84, 	 -75, 	 -73, 	 -67, 	 -68, 	 -63, 	 -62, 	 -62, 	 -57, 	 -56, 	 -52, 	 -45, 	 -43, 	 -41, 	 -37, 	 -40, 	 -53, 	 -53, 	 -40, 	 -30, 	 -38, 	 -41, 	 -43, 	 -43, 	 -31, 	 -24, 	 -34, 	 -74, 	 -79, 	 -81, 	 -82, 	 -83, 	 -85, 	 -86, 	 -86, 	 -88, 	 -89, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 		 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -90, 	 -91, 	 -91, 	 -90, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -92, 	 -92, 	 -91, 	 -91, 	 -92, 	 -90, 	 -90, 	 -85, 	 -71, 	 -60, 	 -39, 	 -15, 	 -18, 	 -26, 	 -67, 	 -62, 	 -14, 	  -7, 	 -16, 	 -58, 	 -83, 	 -88, 	 -76, 	 -38, 	 -62, 	 -68, 	 -53, 	 -70, 	 -60, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -85, 	 -85, 	 -85, 	 -85, 	 -84, 	 -85, 	 -85, 	 -86, 	 -83, 	 -84, 	 -82, 	 -86, 	 -86, 	 -84, 	 -83, 	 -80, 	 -76, 	 -73, 	 -68, 	 -64, 	 -64, 	 -60, 	 -61, 	 -57, 	 -56, 	 -51, 	 -47, 	 -43, 	 -41, 	 -39, 	 -46, 	 -54, 	 -45, 	 -37, 	 -31, 	 -37, 	 -33, 	 -32, 	 -28, 	 -18, 	 -23, 	 -57, 	 -77, 	 -79, 	 -79, 	 -82, 	 -84, 	 -83, 	 -84, 	 -86, 	 -88, 	 -89, 	 -88, 	 -88, 	 -88, 	 -88, 		 -88, 	 -88, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -92, 	 -91, 	 -91, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -88, 	 -90, 	 -91, 	 -91, 	 -91, 	 -91, 	 -92, 	 -92, 	 -93, 	 -92, 	 -92, 	 -91, 	 -87, 	 -75, 	 -63, 	 -46, 	 -16, 	 -23, 	 -29, 	 -45, 	 -38, 	   4, 	   9, 	   9, 	   2, 	 -36, 	 -84, 	 -79, 	 -47, 	 -75, 	 -79, 	 -73, 	 -74, 	 -73, 	
 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -85, 	 -84, 	 -86, 	 -85, 	 -84, 	 -85, 	 -85, 	 -85, 	 -84, 	 -82, 	 -82, 	 -88, 	 -84, 	 -83, 	 -83, 	 -79, 	 -73, 	 -71, 	 -67, 	 -63, 	 -60, 	 -60, 	 -57, 	 -56, 	 -55, 	 -50, 	 -44, 	 -38, 	 -39, 	 -39, 	 -50, 	 -51, 	 -34, 	 -32, 	 -31, 	 -28, 	 -24, 	 -21, 	 -18, 	 -20, 	 -36, 	 -76, 	 -79, 	 -81, 	 -82, 	 -83, 	 -83, 	 -84, 	 -85, 	 -87, 	 -87, 	 -88, 	 -88, 	 -88, 	 -88, 		 -88, 	 -88, 	 -88, 	 -88, 	 -89, 	 -90, 	 -90, 	 -90, 	 -91, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -90, 	 -91, 	 -91, 	 -90, 	 -89, 	 -88, 	 -90, 	 -88, 	 -90, 	 -90, 	 -90, 	 -88, 	 -90, 	 -90, 	 -90, 	 -91, 	 -91, 	 -92, 	 -92, 	 -92, 	 -93, 	 -90, 	 -91, 	 -88, 	 -80, 	 -62, 	 -47, 	 -21, 	 -19, 	 -33, 	 -36, 	 -25, 	  10, 	   6, 	   5, 	   7, 	  -5, 	 -64, 	 -72, 	 -45, 	 -75, 	 -80, 	 -77, 	 -77, 	 -80, 	
 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -83, 	 -84, 	 -84, 	 -85, 	 -85, 	 -85, 	 -85, 	 -82, 	 -83, 	 -85, 	 -84, 	 -82, 	 -83, 	 -76, 	 -71, 	 -69, 	 -65, 	 -64, 	 -61, 	 -60, 	 -60, 	 -58, 	 -53, 	 -49, 	 -44, 	 -39, 	 -39, 	 -46, 	 -51, 	 -43, 	 -29, 	 -23, 	 -24, 	 -19, 	 -21, 	 -20, 	 -18, 	 -30, 	 -60, 	 -76, 	 -79, 	 -80, 	 -81, 	 -82, 	 -83, 	 -85, 	 -85, 	 -86, 	 -87, 	 -87, 	 -87, 	 -87, 		 -87, 	 -87, 	 -87, 	 -88, 	 -89, 	 -88, 	 -88, 	 -89, 	 -90, 	 -90, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -90, 	 -90, 	 -90, 	 -90, 	 -88, 	 -88, 	 -89, 	 -88, 	 -90, 	 -87, 	 -88, 	 -88, 	 -90, 	 -90, 	 -90, 	 -91, 	 -92, 	 -92, 	 -92, 	 -92, 	 -92, 	 -90, 	 -91, 	 -88, 	 -82, 	 -66, 	 -51, 	 -27, 	 -10, 	 -28, 	 -31, 	 -53, 	 -34, 	   1, 	  -4, 	  -6, 	 -18, 	 -72, 	 -74, 	 -46, 	 -72, 	 -72, 	 -61, 	 -28, 	 -66, 	
 -84, 	 -84, 	 -85, 	 -85, 	 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -85, 	 -82, 	 -82, 	 -86, 	 -83, 	 -83, 	 -81, 	 -75, 	 -72, 	 -67, 	 -67, 	 -61, 	 -63, 	 -60, 	 -60, 	 -56, 	 -52, 	 -48, 	 -42, 	 -38, 	 -43, 	 -51, 	 -51, 	 -33, 	 -18, 	 -18, 	 -20, 	 -18, 	 -21, 	 -19, 	 -23, 	 -43, 	 -73, 	 -78, 	 -77, 	 -81, 	 -82, 	 -83, 	 -84, 	 -85, 	 -86, 	 -88, 	 -88, 	 -87, 	 -87, 		 -87, 	 -87, 	 -88, 	 -87, 	 -87, 	 -88, 	 -87, 	 -87, 	 -87, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -88, 	 -90, 	 -89, 	 -89, 	 -88, 	 -89, 	 -88, 	 -90, 	 -86, 	 -90, 	 -86, 	 -86, 	 -88, 	 -89, 	 -89, 	 -90, 	 -91, 	 -92, 	 -91, 	 -94, 	 -93, 	 -90, 	 -91, 	 -90, 	 -89, 	 -82, 	 -70, 	 -54, 	 -31, 	 -12, 	 -18, 	 -14, 	 -55, 	 -74, 	 -70, 	 -59, 	 -53, 	 -66, 	 -83, 	 -79, 	 -59, 	 -73, 	 -69, 	 -68, 	 -28, 	 -36, 	
 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -85, 	 -83, 	 -82, 	 -84, 	 -84, 	 -83, 	 -81, 	 -78, 	 -75, 	 -71, 	 -69, 	 -65, 	 -63, 	 -63, 	 -61, 	 -59, 	 -58, 	 -52, 	 -45, 	 -39, 	 -43, 	 -48, 	 -52, 	 -38, 	 -23, 	 -14, 	 -17, 	 -19, 	 -16, 	 -20, 	 -23, 	 -31, 	 -56, 	 -70, 	 -74, 	 -78, 	 -78, 	 -81, 	 -85, 	 -84, 	 -85, 	 -89, 	 -85, 	 -86, 	 -87, 		 -87, 	 -86, 	 -87, 	 -87, 	 -87, 	 -87, 	 -87, 	 -86, 	 -86, 	 -88, 	 -87, 	 -87, 	 -88, 	 -87, 	 -87, 	 -87, 	 -87, 	 -87, 	 -87, 	 -89, 	 -89, 	 -89, 	 -90, 	 -90, 	 -86, 	 -87, 	 -86, 	 -87, 	 -85, 	 -87, 	 -86, 	 -85, 	 -89, 	 -89, 	 -92, 	 -91, 	 -92, 	 -92, 	 -91, 	 -87, 	 -89, 	 -88, 	 -89, 	 -88, 	 -73, 	 -59, 	 -38, 	 -11, 	 -10, 	  -8, 	 -33, 	 -82, 	 -83, 	 -83, 	 -83, 	 -84, 	 -87, 	 -74, 	 -46, 	 -59, 	 -71, 	 -68, 	 -58, 	 -59, 	
 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -84, 	 -83, 	 -83, 	 -83, 	 -83, 	 -84, 	 -84, 	 -84, 	 -85, 	 -84, 	 -82, 	 -82, 	 -85, 	 -83, 	 -82, 	 -79, 	 -76, 	 -72, 	 -69, 	 -69, 	 -64, 	 -64, 	 -61, 	 -60, 	 -61, 	 -56, 	 -47, 	 -41, 	 -42, 	 -46, 	 -51, 	 -45, 	 -31, 	 -13, 	 -20, 	 -17, 	 -20, 	 -20, 	 -17, 	 -28, 	 -41, 	 -62, 	 -63, 	 -68, 	 -73, 	 -76, 	 -81, 	 -84, 	 -85, 	 -85, 	 -84, 	 -86, 	 -86, 		 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -87, 	 -86, 	 -87, 	 -87, 	 -86, 	 -86, 	 -87, 	 -86, 	 -85, 	 -81, 	 -82, 	 -85, 	 -82, 	 -83, 	 -83, 	 -85, 	 -88, 	 -89, 	 -89, 	 -93, 	 -91, 	 -90, 	 -88, 	 -86, 	 -87, 	 -89, 	 -89, 	 -84, 	 -78, 	 -61, 	 -46, 	 -28, 	 -18, 	 -28, 	 -15, 	 -75, 	 -81, 	 -83, 	 -85, 	 -61, 	 -20, 	  -2, 	  13, 	  15, 	  20, 	  31, 	  14, 	 -45, 	
 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -83, 	 -82, 	 -82, 	 -82, 	 -83, 	 -83, 	 -82, 	 -83, 	 -83, 	 -83, 	 -84, 	 -84, 	 -86, 	 -81, 	 -83, 	 -83, 	 -86, 	 -81, 	 -84, 	 -80, 	 -76, 	 -72, 	 -68, 	 -69, 	 -66, 	 -62, 	 -62, 	 -60, 	 -59, 	 -49, 	 -42, 	 -45, 	 -44, 	 -49, 	 -50, 	 -36, 	 -16, 	 -14, 	 -18, 	 -15, 	 -17, 	 -18, 	 -18, 	 -29, 	 -48, 	 -57, 	 -66, 	 -66, 	 -69, 	 -73, 	 -81, 	 -85, 	 -85, 	 -87, 	 -87, 	 -85, 		 -87, 	 -86, 	 -85, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -86, 	 -85, 	 -85, 	 -85, 	 -85, 	 -86, 	 -84, 	 -86, 	 -85, 	 -83, 	 -87, 	 -82, 	 -81, 	 -80, 	 -73, 	 -56, 	 -53, 	 -55, 	 -61, 	 -62, 	 -65, 	 -68, 	 -76, 	 -64, 	 -73, 	 -90, 	 -92, 	 -91, 	 -90, 	 -89, 	 -89, 	 -92, 	 -90, 	 -88, 	 -78, 	 -60, 	 -47, 	 -31, 	 -25, 	 -36, 	  -7, 	 -27, 	 -46, 	 -40, 	 -42, 	 -24, 	  -5, 	  -1, 	 -31, 	 -24, 	  12, 	  39, 	  15, 	 -29, 	
 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -83, 	 -82, 	 -83, 	 -81, 	 -82, 	 -83, 	 -85, 	 -84, 	 -83, 	 -84, 	 -84, 	 -83, 	 -81, 	 -86, 	 -85, 	 -82, 	 -81, 	 -76, 	 -75, 	 -69, 	 -67, 	 -64, 	 -66, 	 -61, 	 -60, 	 -60, 	 -51, 	 -44, 	 -45, 	 -47, 	 -48, 	 -48, 	 -42, 	 -25, 	 -15, 	 -13, 	 -15, 	 -18, 	 -24, 	 -22, 	 -25, 	 -38, 	 -54, 	 -58, 	 -63, 	 -62, 	 -57, 	 -71, 	 -77, 	 -82, 	 -85, 	 -84, 	 -85, 		 -85, 	 -86, 	 -86, 	 -85, 	 -86, 	 -85, 	 -84, 	 -85, 	 -87, 	 -87, 	 -86, 	 -84, 	 -82, 	 -84, 	 -85, 	 -85, 	 -84, 	 -82, 	 -79, 	 -80, 	 -82, 	 -85, 	 -84, 	 -82, 	 -73, 	 -58, 	 -47, 	 -50, 	 -53, 	 -56, 	 -56, 	 -55, 	 -61, 	 -55, 	 -70, 	 -88, 	 -93, 	 -89, 	 -89, 	 -87, 	 -89, 	 -93, 	 -89, 	 -91, 	 -86, 	 -67, 	 -49, 	 -34, 	 -28, 	 -39, 	 -15, 	 -25, 	 -34, 	 -31, 	 -25, 	 -31, 	   5, 	  27, 	  13, 	  -4, 	 -22, 	  10, 	  26, 	  20, 	
 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -83, 	 -82, 	 -81, 	 -81, 	 -82, 	 -82, 	 -81, 	 -82, 	 -84, 	 -83, 	 -83, 	 -83, 	 -81, 	 -84, 	 -84, 	 -83, 	 -84, 	 -79, 	 -77, 	 -71, 	 -68, 	 -67, 	 -65, 	 -65, 	 -61, 	 -63, 	 -54, 	 -47, 	 -42, 	 -47, 	 -46, 	 -47, 	 -48, 	 -32, 	  -9, 	 -16, 	 -18, 	 -23, 	 -26, 	 -27, 	 -29, 	 -34, 	 -45, 	 -53, 	 -57, 	 -60, 	 -51, 	 -56, 	 -58, 	 -63, 	 -71, 	 -77, 	 -82, 		 -83, 	 -84, 	 -85, 	 -84, 	 -84, 	 -83, 	 -84, 	 -84, 	 -84, 	 -85, 	 -86, 	 -85, 	 -83, 	 -85, 	 -83, 	 -81, 	 -80, 	 -76, 	 -75, 	 -72, 	 -74, 	 -80, 	 -85, 	 -82, 	 -78, 	 -67, 	 -54, 	 -59, 	 -53, 	 -56, 	 -53, 	 -54, 	 -53, 	 -49, 	 -57, 	 -81, 	 -90, 	 -86, 	 -87, 	 -88, 	 -89, 	 -90, 	 -91, 	 -91, 	 -87, 	 -71, 	 -46, 	 -36, 	 -31, 	 -34, 	 -16, 	 -24, 	 -70, 	 -66, 	 -62, 	 -41, 	  -5, 	  16, 	  35, 	  26, 	  34, 	  38, 	  35, 	  41, 	
 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -83, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -81, 	 -81, 	 -80, 	 -80, 	 -80, 	 -81, 	 -82, 	 -82, 	 -83, 	 -83, 	 -82, 	 -83, 	 -81, 	 -85, 	 -83, 	 -83, 	 -80, 	 -75, 	 -72, 	 -68, 	 -67, 	 -65, 	 -65, 	 -61, 	 -64, 	 -55, 	 -47, 	 -39, 	 -44, 	 -42, 	 -45, 	 -50, 	 -40, 	 -18, 	 -19, 	 -25, 	 -27, 	 -27, 	 -30, 	 -31, 	 -36, 	 -41, 	 -50, 	 -54, 	 -54, 	 -50, 	 -50, 	 -55, 	 -59, 	 -58, 	 -61, 	 -71, 		 -77, 	 -78, 	 -80, 	 -84, 	 -84, 	 -83, 	 -83, 	 -84, 	 -85, 	 -83, 	 -84, 	 -83, 	 -79, 	 -79, 	 -73, 	 -70, 	 -73, 	 -71, 	 -71, 	 -72, 	 -70, 	 -77, 	 -82, 	 -82, 	 -77, 	 -70, 	 -64, 	 -65, 	 -60, 	 -56, 	 -51, 	 -49, 	 -45, 	 -48, 	 -54, 	 -73, 	 -81, 	 -85, 	 -85, 	 -86, 	 -90, 	 -91, 	 -90, 	 -91, 	 -87, 	 -78, 	 -42, 	 -41, 	 -46, 	 -29, 	 -30, 	 -26, 	 -70, 	 -80, 	 -61, 	 -50, 	 -50, 	 -26, 	  12, 	  11, 	  33, 	  26, 	 -25, 	  37, 	
 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -81, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -80, 	 -80, 	 -80, 	 -80, 	 -79, 	 -80, 	 -81, 	 -81, 	 -82, 	 -83, 	 -81, 	 -83, 	 -81, 	 -85, 	 -86, 	 -83, 	 -81, 	 -78, 	 -74, 	 -70, 	 -70, 	 -66, 	 -65, 	 -63, 	 -64, 	 -56, 	 -44, 	 -35, 	 -38, 	 -40, 	 -43, 	 -50, 	 -43, 	 -29, 	 -22, 	 -29, 	 -30, 	 -30, 	 -32, 	 -36, 	 -42, 	 -46, 	 -46, 	 -49, 	 -53, 	 -46, 	 -51, 	 -54, 	 -62, 	 -63, 	 -67, 	 -75, 		 -77, 	 -78, 	 -81, 	 -83, 	 -82, 	 -83, 	 -83, 	 -82, 	 -83, 	 -82, 	 -83, 	 -80, 	 -72, 	 -69, 	 -58, 	 -56, 	 -59, 	 -59, 	 -61, 	 -66, 	 -58, 	 -61, 	 -67, 	 -70, 	 -72, 	 -70, 	 -63, 	 -64, 	 -64, 	 -66, 	 -57, 	 -51, 	 -45, 	 -42, 	 -36, 	 -66, 	 -72, 	 -73, 	 -81, 	 -87, 	 -89, 	 -91, 	 -90, 	 -90, 	 -87, 	 -82, 	 -49, 	 -31, 	 -42, 	 -34, 	 -29, 	 -23, 	 -52, 	 -64, 	 -57, 	 -63, 	 -66, 	 -71, 	 -69, 	 -37, 	 -22, 	   1, 	 -28, 	  -7, 	
 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -82, 	 -83, 	 -81, 	 -81, 	 -81, 	 -80, 	 -79, 	 -79, 	 -79, 	 -79, 	 -79, 	 -78, 	 -78, 	 -79, 	 -81, 	 -81, 	 -82, 	 -83, 	 -83, 	 -83, 	 -85, 	 -85, 	 -81, 	 -80, 	 -72, 	 -70, 	 -68, 	 -65, 	 -65, 	 -63, 	 -63, 	 -57, 	 -44, 	 -33, 	 -34, 	 -35, 	 -43, 	 -45, 	 -47, 	 -35, 	 -26, 	 -31, 	 -31, 	 -31, 	 -33, 	 -37, 	 -43, 	 -49, 	 -52, 	 -57, 	 -61, 	 -54, 	 -57, 	 -61, 	 -65, 	 -66, 	 -71, 	 -73, 		 -79, 	 -79, 	 -81, 	 -83, 	 -82, 	 -79, 	 -83, 	 -79, 	 -78, 	 -78, 	 -62, 	 -56, 	 -44, 	 -38, 	 -29, 	 -35, 	 -40, 	 -46, 	 -47, 	 -51, 	 -54, 	 -47, 	 -53, 	 -59, 	 -64, 	 -70, 	 -66, 	 -68, 	 -65, 	 -71, 	 -65, 	 -56, 	 -52, 	 -46, 	 -30, 	 -57, 	 -64, 	 -65, 	 -74, 	 -87, 	 -89, 	 -90, 	 -91, 	 -90, 	 -86, 	 -80, 	 -64, 	 -41, 	 -47, 	 -45, 	 -37, 	 -36, 	 -40, 	 -41, 	 -45, 	 -40, 	 -49, 	 -61, 	 -85, 	 -75, 	 -71, 	 -47, 	 -33, 	 -49, 	
 -81, 	 -81, 	 -81, 	 -81, 	 -81, 	 -81, 	 -81, 	 -82, 	 -81, 	 -81, 	 -81, 	 -80, 	 -79, 	 -79, 	 -79, 	 -79, 	 -78, 	 -77, 	 -78, 	 -78, 	 -78, 	 -79, 	 -81, 	 -81, 	 -82, 	 -82, 	 -82, 	 -84, 	 -82, 	 -80, 	 -75, 	 -70, 	 -68, 	 -65, 	 -64, 	 -62, 	 -63, 	 -59, 	 -49, 	 -34, 	 -31, 	 -34, 	 -38, 	 -44, 	 -51, 	 -42, 	 -31, 	 -29, 	 -35, 	 -31, 	 -34, 	 -41, 	 -48, 	 -52, 	 -60, 	 -61, 	 -65, 	 -60, 	 -53, 	 -58, 	 -64, 	 -68, 	 -67, 	 -69, 		 -74, 	 -72, 	 -70, 	 -69, 	 -64, 	 -62, 	 -57, 	 -52, 	 -52, 	 -37, 	 -31, 	 -31, 	 -27, 	 -27, 	 -23, 	 -31, 	 -37, 	 -42, 	 -48, 	 -50, 	 -52, 	 -42, 	 -49, 	 -50, 	 -55, 	 -61, 	 -65, 	 -64, 	 -70, 	 -68, 	 -71, 	 -63, 	 -44, 	 -29, 	 -18, 	 -36, 	 -41, 	 -39, 	 -45, 	 -48, 	 -54, 	 -66, 	 -82, 	 -88, 	 -87, 	 -84, 	 -74, 	 -56, 	 -58, 	 -60, 	 -61, 	 -61, 	 -61, 	 -50, 	 -62, 	 -56, 	 -49, 	 -63, 	 -85, 	 -86, 	 -84, 	 -81, 	 -73, 	 -70, 	
 -81, 	 -81, 	 -81, 	 -82, 	 -81, 	 -81, 	 -82, 	 -82, 	 -81, 	 -81, 	 -81, 	 -80, 	 -79, 	 -79, 	 -79, 	 -79, 	 -78, 	 -77, 	 -77, 	 -78, 	 -77, 	 -76, 	 -79, 	 -79, 	 -81, 	 -83, 	 -81, 	 -84, 	 -83, 	 -81, 	 -79, 	 -70, 	 -66, 	 -65, 	 -63, 	 -61, 	 -62, 	 -61, 	 -50, 	 -39, 	 -32, 	 -29, 	 -36, 	 -41, 	 -47, 	 -44, 	 -40, 	 -34, 	 -37, 	 -35, 	 -42, 	 -48, 	 -53, 	 -65, 	 -68, 	 -68, 	 -69, 	 -67, 	 -56, 	 -58, 	 -57, 	 -56, 	 -51, 	 -49, 		 -41, 	 -38, 	 -28, 	 -24, 	 -21, 	 -21, 	 -21, 	 -20, 	 -23, 	 -24, 	 -23, 	 -28, 	 -26, 	 -25, 	 -26, 	 -27, 	 -39, 	 -44, 	 -54, 	 -52, 	 -54, 	 -41, 	 -44, 	 -47, 	 -48, 	 -53, 	 -62, 	 -65, 	 -66, 	 -72, 	 -73, 	 -66, 	 -48, 	 -43, 	 -50, 	 -50, 	 -58, 	 -49, 	 -55, 	 -47, 	 -48, 	 -54, 	 -75, 	 -87, 	 -86, 	 -84, 	 -78, 	 -69, 	 -64, 	 -78, 	 -61, 	 -47, 	 -69, 	 -72, 	 -66, 	 -64, 	 -67, 	 -84, 	 -88, 	 -85, 	 -85, 	 -72, 	 -66, 	 -62, 	
 -81, 	 -82, 	 -82, 	 -82, 	 -83, 	 -82, 	 -83, 	 -82, 	 -84, 	 -83, 	 -82, 	 -83, 	 -82, 	 -81, 	 -80, 	 -80, 	 -78, 	 -78, 	 -79, 	 -79, 	 -80, 	 -78, 	 -79, 	 -79, 	 -80, 	 -81, 	 -83, 	 -81, 	 -86, 	 -80, 	 -80, 	 -73, 	 -67, 	 -65, 	 -65, 	 -65, 	 -60, 	 -58, 	 -56, 	 -44, 	 -31, 	 -29, 	 -31, 	 -41, 	 -45, 	 -49, 	 -42, 	 -40, 	 -39, 	 -36, 	 -43, 	 -53, 	 -60, 	 -65, 	 -70, 	 -70, 	 -73, 	 -66, 	 -57, 	 -56, 	 -55, 	 -52, 	 -50, 	 -45, 		 -37, 	 -31, 	 -18, 	 -22, 	 -21, 	 -14, 	 -17, 	 -17, 	 -23, 	 -22, 	 -21, 	 -23, 	 -29, 	 -28, 	 -29, 	 -32, 	 -41, 	 -52, 	 -56, 	 -57, 	 -59, 	 -47, 	 -37, 	 -44, 	 -42, 	 -46, 	 -52, 	 -57, 	 -64, 	 -68, 	 -72, 	 -71, 	 -68, 	 -72, 	 -72, 	 -67, 	 -65, 	 -70, 	 -69, 	 -67, 	 -68, 	 -72, 	 -85, 	 -81, 	 -74, 	 -67, 	 -53, 	 -69, 	 -71, 	 -76, 	 -71, 	 -45, 	 -62, 	 -64, 	 -56, 	 -51, 	 -60, 	 -83, 	 -87, 	 -88, 	 -77, 	 -57, 	 -61, 	 -53, 	
 -81, 	 -82, 	 -82, 	 -83, 	 -84, 	 -83, 	 -83, 	 -82, 	 -82, 	 -83, 	 -83, 	 -83, 	 -82, 	 -82, 	 -81, 	 -79, 	 -79, 	 -80, 	 -78, 	 -78, 	 -78, 	 -77, 	 -78, 	 -78, 	 -79, 	 -79, 	 -82, 	 -80, 	 -84, 	 -82, 	 -80, 	 -74, 	 -70, 	 -65, 	 -64, 	 -64, 	 -60, 	 -59, 	 -54, 	 -46, 	 -33, 	 -30, 	 -31, 	 -38, 	 -44, 	 -50, 	 -42, 	 -42, 	 -37, 	 -40, 	 -44, 	 -53, 	 -63, 	 -64, 	 -74, 	 -71, 	 -72, 	 -65, 	 -55, 	 -53, 	 -52, 	 -50, 	 -50, 	 -42, 		 -33, 	 -24, 	 -26, 	 -16, 	 -19, 	 -12, 	 -20, 	 -13, 	 -21, 	 -20, 	 -18, 	 -24, 	 -32, 	 -31, 	 -29, 	 -36, 	 -45, 	 -57, 	 -56, 	 -60, 	 -58, 	 -50, 	 -35, 	 -37, 	 -37, 	 -40, 	 -40, 	 -49, 	 -54, 	 -66, 	 -69, 	 -72, 	 -79, 	 -78, 	 -84, 	 -69, 	 -72, 	 -75, 	 -66, 	 -56, 	 -56, 	 -70, 	 -83, 	 -67, 	 -29, 	 -40, 	 -59, 	 -79, 	 -67, 	 -62, 	 -77, 	 -53, 	 -57, 	 -58, 	 -55, 	 -51, 	 -58, 	 -83, 	 -85, 	 -88, 	 -81, 	 -70, 	 -76, 	 -72, 	
 -82, 	 -82, 	 -82, 	 -84, 	 -83, 	 -83, 	 -84, 	 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -82, 	 -82, 	 -79, 	 -80, 	 -78, 	 -79, 	 -78, 	 -79, 	 -78, 	 -78, 	 -78, 	 -82, 	 -80, 	 -84, 	 -84, 	 -82, 	 -79, 	 -72, 	 -65, 	 -65, 	 -62, 	 -60, 	 -57, 	 -56, 	 -48, 	 -41, 	 -33, 	 -29, 	 -36, 	 -41, 	 -51, 	 -46, 	 -43, 	 -39, 	 -40, 	 -43, 	 -56, 	 -64, 	 -71, 	 -74, 	 -72, 	 -70, 	 -63, 	 -52, 	 -50, 	 -47, 	 -44, 	 -45, 	 -38, 		 -29, 	 -25, 	 -25, 	 -19, 	 -21, 	 -13, 	 -20, 	 -19, 	 -18, 	 -19, 	 -15, 	 -26, 	 -27, 	 -36, 	 -29, 	 -39, 	 -45, 	 -54, 	 -57, 	 -66, 	 -63, 	 -52, 	 -39, 	 -38, 	 -35, 	 -34, 	 -39, 	 -41, 	 -46, 	 -60, 	 -62, 	 -71, 	 -75, 	 -82, 	 -80, 	 -77, 	 -71, 	 -67, 	 -53, 	 -45, 	 -47, 	 -60, 	 -66, 	 -64, 	 -57, 	 -42, 	 -73, 	 -85, 	 -39, 	 -47, 	 -78, 	 -71, 	 -57, 	 -59, 	 -57, 	 -54, 	 -58, 	 -71, 	 -88, 	 -85, 	 -78, 	 -73, 	 -72, 	 -63, 	
 -82, 	 -83, 	 -83, 	 -84, 	 -83, 	 -84, 	 -84, 	 -82, 	 -82, 	 -84, 	 -83, 	 -84, 	 -84, 	 -83, 	 -83, 	 -83, 	 -84, 	 -81, 	 -81, 	 -80, 	 -80, 	 -81, 	 -80, 	 -79, 	 -79, 	 -81, 	 -80, 	 -81, 	 -82, 	 -84, 	 -82, 	 -80, 	 -73, 	 -66, 	 -65, 	 -62, 	 -60, 	 -57, 	 -56, 	 -52, 	 -44, 	 -35, 	 -30, 	 -33, 	 -41, 	 -52, 	 -49, 	 -44, 	 -41, 	 -47, 	 -49, 	 -59, 	 -67, 	 -74, 	 -73, 	 -71, 	 -68, 	 -60, 	 -49, 	 -45, 	 -40, 	 -40, 	 -42, 	 -34, 		 -27, 	 -26, 	 -25, 	 -23, 	 -16, 	 -17, 	 -17, 	 -19, 	 -19, 	 -17, 	 -16, 	 -24, 	 -28, 	 -35, 	 -31, 	 -43, 	 -44, 	 -56, 	 -57, 	 -64, 	 -62, 	 -58, 	 -38, 	 -35, 	 -33, 	 -34, 	 -32, 	 -36, 	 -42, 	 -48, 	 -55, 	 -61, 	 -64, 	 -52, 	 -65, 	 -80, 	 -74, 	 -61, 	 -45, 	 -26, 	 -36, 	 -52, 	 -47, 	 -14, 	 -34, 	 -32, 	 -41, 	 -68, 	 -24, 	 -60, 	 -69, 	 -82, 	 -64, 	 -62, 	 -55, 	 -53, 	 -48, 	 -57, 	 -83, 	 -72, 	 -50, 	 -62, 	 -55, 	 -30, 	
 -82, 	 -82, 	 -82, 	 -82, 	 -84, 	 -82, 	 -84, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -82, 	 -81, 	 -80, 	 -81, 	 -80, 	 -81, 	 -80, 	 -78, 	 -79, 	 -78, 	 -82, 	 -84, 	 -80, 	 -73, 	 -68, 	 -66, 	 -63, 	 -61, 	 -59, 	 -55, 	 -52, 	 -48, 	 -38, 	 -36, 	 -33, 	 -35, 	 -48, 	 -53, 	 -43, 	 -40, 	 -45, 	 -53, 	 -60, 	 -68, 	 -73, 	 -75, 	 -67, 	 -62, 	 -56, 	 -49, 	 -39, 	 -33, 	 -31, 	 -33, 	 -31, 		 -32, 	 -26, 	 -22, 	 -23, 	 -19, 	 -18, 	 -15, 	 -19, 	 -17, 	 -18, 	 -18, 	 -25, 	 -26, 	 -35, 	 -35, 	 -41, 	 -46, 	 -56, 	 -60, 	 -65, 	 -63, 	 -55, 	 -39, 	 -35, 	 -34, 	 -30, 	 -28, 	 -34, 	 -35, 	 -44, 	 -50, 	 -59, 	 -47, 	 -12, 	 -71, 	 -82, 	 -79, 	 -62, 	 -50, 	 -22, 	 -32, 	 -46, 	 -50, 	 -34, 	 -28, 	 -37, 	 -33, 	 -44, 	 -45, 	 -53, 	 -60, 	 -80, 	 -62, 	 -62, 	 -56, 	 -52, 	 -51, 	 -57, 	 -71, 	 -68, 	 -59, 	 -59, 	 -59, 	 -52, 	
 -82, 	 -83, 	 -82, 	 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -81, 	 -82, 	 -83, 	 -81, 	 -82, 	 -82, 	 -82, 	 -81, 	 -80, 	 -80, 	 -80, 	 -80, 	 -84, 	 -81, 	 -79, 	 -72, 	 -65, 	 -64, 	 -62, 	 -61, 	 -59, 	 -53, 	 -50, 	 -43, 	 -37, 	 -34, 	 -36, 	 -44, 	 -51, 	 -46, 	 -43, 	 -44, 	 -52, 	 -59, 	 -67, 	 -66, 	 -67, 	 -61, 	 -57, 	 -50, 	 -42, 	 -35, 	 -27, 	 -27, 	 -33, 	 -31, 		 -30, 	 -27, 	 -21, 	 -23, 	 -19, 	 -18, 	 -20, 	 -19, 	 -20, 	 -20, 	 -21, 	 -26, 	 -24, 	 -35, 	 -37, 	 -41, 	 -47, 	 -57, 	 -66, 	 -64, 	 -61, 	 -56, 	 -39, 	 -33, 	 -36, 	 -33, 	 -30, 	 -31, 	 -32, 	 -40, 	 -42, 	 -49, 	 -42, 	 -44, 	 -72, 	 -82, 	 -82, 	 -64, 	 -58, 	 -39, 	 -40, 	 -47, 	 -60, 	 -64, 	 -46, 	 -43, 	 -22, 	 -40, 	 -67, 	 -56, 	 -58, 	 -78, 	 -63, 	 -61, 	 -57, 	 -49, 	 -51, 	 -52, 	 -54, 	 -63, 	 -62, 	 -64, 	 -55, 	 -59, 	
 -81, 	 -83, 	 -82, 	 -82, 	 -83, 	 -83, 	 -83, 	 -84, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -84, 	 -83, 	 -83, 	 -84, 	 -83, 	 -82, 	 -83, 	 -82, 	 -84, 	 -84, 	 -82, 	 -80, 	 -80, 	 -79, 	 -84, 	 -84, 	 -81, 	 -74, 	 -67, 	 -67, 	 -64, 	 -61, 	 -61, 	 -54, 	 -51, 	 -46, 	 -40, 	 -38, 	 -36, 	 -42, 	 -53, 	 -49, 	 -39, 	 -37, 	 -49, 	 -54, 	 -65, 	 -63, 	 -65, 	 -58, 	 -51, 	 -45, 	 -37, 	 -32, 	 -24, 	 -27, 	 -32, 	 -32, 		 -32, 	 -28, 	 -26, 	 -21, 	 -22, 	 -20, 	 -18, 	 -21, 	 -21, 	 -20, 	 -25, 	 -25, 	 -23, 	 -30, 	 -43, 	 -46, 	 -50, 	 -61, 	 -65, 	 -64, 	 -61, 	 -50, 	 -43, 	 -30, 	 -38, 	 -37, 	 -34, 	 -31, 	 -29, 	 -35, 	 -36, 	 -41, 	 -46, 	 -51, 	 -71, 	 -76, 	 -78, 	 -62, 	 -58, 	 -44, 	 -46, 	 -49, 	 -61, 	 -75, 	 -67, 	 -43, 	 -35, 	 -23, 	 -32, 	 -50, 	 -35, 	 -64, 	 -69, 	 -61, 	 -57, 	 -50, 	 -52, 	 -50, 	 -53, 	 -71, 	 -71, 	 -61, 	 -59, 	 -62, 	
 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -81, 	 -80, 	 -79, 	 -81, 	 -84, 	 -80, 	 -76, 	 -72, 	 -67, 	 -66, 	 -64, 	 -62, 	 -57, 	 -55, 	 -53, 	 -41, 	 -44, 	 -38, 	 -47, 	 -53, 	 -53, 	 -39, 	 -33, 	 -44, 	 -51, 	 -59, 	 -58, 	 -56, 	 -53, 	 -44, 	 -37, 	 -27, 	 -23, 	 -21, 	 -25, 	 -30, 	 -31, 		 -31, 	 -25, 	 -24, 	 -24, 	 -25, 	 -15, 	 -19, 	 -20, 	 -23, 	 -26, 	 -27, 	 -16, 	 -20, 	 -34, 	 -44, 	 -46, 	 -59, 	 -59, 	 -66, 	 -63, 	 -59, 	 -54, 	 -44, 	 -34, 	 -37, 	 -38, 	 -32, 	 -29, 	 -36, 	 -32, 	 -32, 	 -37, 	 -46, 	 -53, 	 -67, 	 -70, 	 -74, 	 -65, 	 -61, 	 -47, 	 -45, 	 -46, 	 -65, 	 -80, 	 -80, 	 -58, 	 -64, 	 -63, 	 -50, 	 -42, 	 -44, 	 -59, 	 -73, 	 -59, 	 -56, 	 -49, 	 -47, 	 -49, 	 -58, 	 -67, 	 -73, 	 -66, 	 -64, 	 -65, 	
 -82, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -82, 	 -82, 	 -83, 	 -83, 	 -83, 	 -84, 	 -84, 	 -84, 	 -84, 	 -84, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -83, 	 -82, 	 -83, 	 -79, 	 -78, 	 -78, 	 -85, 	 -81, 	 -79, 	 -73, 	 -67, 	 -66, 	 -64, 	 -62, 	 -60, 	 -58, 	 -55, 	 -45, 	 -44, 	 -38, 	 -42, 	 -51, 	 -56, 	 -39, 	 -32, 	 -34, 	 -46, 	 -52, 	 -50, 	 -51, 	 -47, 	 -40, 	 -31, 	 -24, 	 -21, 	 -21, 	 -26, 	 -30, 	 -31, 		 -28, 	 -29, 	 -21, 	 -17, 	 -23, 	 -15, 	 -21, 	 -19, 	 -26, 	 -29, 	 -29, 	 -18, 	 -20, 	 -37, 	 -49, 	 -52, 	 -63, 	 -63, 	 -66, 	 -65, 	 -60, 	 -57, 	 -46, 	 -38, 	 -38, 	 -43, 	 -33, 	 -33, 	 -32, 	 -32, 	 -33, 	 -39, 	 -42, 	 -40, 	 -34, 	 -31, 	 -54, 	 -63, 	 -60, 	 -49, 	 -46, 	 -49, 	 -71, 	 -75, 	 -83, 	 -79, 	 -78, 	 -64, 	 -50, 	 -35, 	 -35, 	 -59, 	 -73, 	 -61, 	 -52, 	 -48, 	 -48, 	 -46, 	 -47, 	 -71, 	 -71, 	 -66, 	 -63, 	 -65

 };
	
	wire	[7:0] 	row = aa /`TILE_WIDTH;
	wire	[7:0] 	col = aa % `TILE_WIDTH;
	always @(`CLK_RST_EDGE)
		if (`RST)	qa <= 0;
		else if (!cena)		qa <= { mem[row *2*`TILE_WIDTH + col][`W1:0], mem[row *2*`TILE_WIDTH + col + `TILE_WIDTH ][`W1:0]};
endmodule



module coeff_rom(
	input			clk,
	input			rstn,
	input	[13:0]	aa,
	input			cena,
	output reg		[`W_WT1P*4-1:0]	qa
	);

	logic [0:`TILE_WIDTH*`TILE_WIDTH-1][31:0] mem	 = {
 256,	-896,	-4096,	-640,	 832,	3200,	3328,	-1344,	
 576,	2624,	1600,	-2752,	4416,	-1408,	2176,	-3584,	
   0,	 832,	 256,	-5504,	6720,	-9344,	-1984,	-1792,	
-2560,	2432,	6144,	1344,	-960,	5184,	1472,	1024,	
-2880,	1600,	-1024,	-1280,	3008,	-2304,	-960,	-1984,	
4672,	 320,	5504,	 704,	-3904,	4800,	1792,	-448,	
-4160,	-1856,	-2048,	-512,	 256,	-3520,	-3392,	1408,	
-2176,	  64,	1280,	1920,	-3392,	-2752,	-1408,	-1728,

1984,	5760,	5760,	-2304,	1600,	-1728,	-1920,	3456,	
-7104,	-3968,	-2688,	1728,	1856,	 128,	5632,	-1920,	
-2176,	-6208,	 448,	 384,	-2240,	3392,	-3648,	-9024,	
7104,	6528,	2560,	6592,	-832,	-4672,	-4224,	7552,	
-12416,	 320,	-1088,	-3904,	6272,	7744,	4800,	6464,	
1792,	 256,	-4224,	-896,	4480,	1344,	7040,	-5696,	
2560,	-960,	2112,	1088,	2304,	-1280,	 832,	-704,	
-9152,	-4800,	-4928,	2304,	-704,	7936,	1408,	2688,

11072,	3520,	-5440,	3904,	-7616,	3264,	4032,	-7296,	
2368,	-8768,	-3136,	10112,	-4096,	 192,	3840,	2048,	
2560,	-7168,	2048,	 384,	5888,	-5312,	7552,	4736,	
-4032,	-5504,	-6592,	-4736,	8896,	3840,	-5824,	2240,	
-1472,	-192,	-320,	 896,	1728,	-4608,	-1856,	4288,	
1024,	-1792,	4992,	-7552,	-2752,	-6464,	-4288,	1664,	
2304,	-2368,	-4992,	-6912,	4992,	9536,	-4352,	7360,	
-4160,	-2240,	-512,	-11200,	 256,	2048,	-3264,	6912,

7488,	-8064,	-512,	-1280,	1920,	-6528,	-5248,	-640,	
-5184,	 448,	12992,	 192,	-4224,	  64,	-10624,	-3776,	
9920,	4736,	3456,	-7360,	2752,	6016,	-256,	-9536,	
 768,	14144,	2176,	2880,	-4288,	13056,	-5952,	-2944,	
1984,	9280,	11904,	-1856,	-11584,	6272,	-2688,	-13760,	
14464,	8704,	13504,	3968,	-960,	9664,	 832,	-12928,	
9600,	2816,	8384,	-7552,	-7232,	8832,	-4352,	-13888,	
6784,	14144,	10048,	3136,	4544,	2688,	13888,	3776

	};

	logic [0:3][0:`TILE_WIDTH/2/4-1][0:`TILE_WIDTH/2-1][0:3][`W_WT1P-1:0] coeff_mem;
	logic	[0:`TILE_WIDTH*`TILE_WIDTH/4-1][`W_WT1P*4-1:0] coeff_mem_4x;
	assign	coeff_mem_4x = coeff_mem;
	initial begin
		for(int cb=0; cb < 4; cb=cb+1) begin
			for(int h = 0; h < `TILE_WIDTH/2/4; h=h+1) begin
				for(int w = 0; w < `TILE_WIDTH/2; w=w+1) begin
					coeff_mem[cb][h][w][0] = 	mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 0 ) + w][31] ? (0 -  mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 0 ) + w] /64) | 1<<`W_WT1 : mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 0 ) + w] /64; 
					coeff_mem[cb][h][w][1] = 	mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 1 ) + w][31] ? (0 -  mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 1 ) + w] /64) | 1<<`W_WT1 : mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 1 ) + w] /64; 
					coeff_mem[cb][h][w][2] = 	mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 2 ) + w][31] ? (0 -  mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 2 ) + w] /64) | 1<<`W_WT1 : mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 2 ) + w] /64; 
					coeff_mem[cb][h][w][3] = 	mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 3 ) + w][31] ? (0 -  mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 3 ) + w] /64) | 1<<`W_WT1 : mem[ cb*(`TILE_WIDTH*`TILE_WIDTH)/4 +  (`TILE_WIDTH/2)*(h*4 + 3 ) + w] /64; 
						
			
								
				end 
			end
		end
	end

	always @(`CLK_RST_EDGE)
		if (`RST)	qa <= 0;
		else if (!cena)		qa <= coeff_mem_4x[aa];
endmodule
interface itf(input clk);
	logic					first_row;
	logic					second_row;
	logic					last_row;
	logic					one_plus_row;
	logic					row_start	;
	logic					row_end	;
	logic					en		;	
	logic		[`W_WT1:0]		x0;
	logic		[`W_WT1:0]		x1;
	logic		[`W_WT1:0]		x2;
	logic		[`W_WT1:0]		x3;
	logic					go;

	logic					plane_start;
	logic					plane_end;
	logic		[3:0]		bit_pos;
	logic 					mq_ready;
	
	
	clocking cb@( `CLK_EDGE);
		output	en;
		//input 	ready;
	endclocking	
	task init();
		en		 <= 0;
		go 		<= 0;
		x0 <= 0;
		x1 <= 0;
		x2 <= 0;
		x3 <= 0;
		first_row <= 0;
		second_row <= 0;
		row_start <= 0;
		row_end	<= 0;
		plane_start <= 0;
		plane_end <= 0;
		bit_pos <= 0;
	endtask
	task drive();
		@cb;
		@cb;
		@cb;
		go <= 1;
		@cb;
		go <= 0;
		@cb;
	endtask
	
	//task drive_frame(logic [`MAX_PATH*8-1:0]	sequence_name; , int nframe);
	
	task start();

		// `define CB_WIDTH 64
		// `define CB_WIDTH 16
		`define CB_WIDTH 8
		// `define CB_WIDTH 4
		// `define START_POS 7
		`define START_POS 7

		logic [0:`CB_WIDTH-1][0:`CB_WIDTH-1][31:0] src = {
11072,	3520,	-5440,	3904,	-7616,	3264,	4032,	-7296,	
2368,	-8768,	-3136,	10112,	-4096,	 192,	3840,	2048,	
2560,	-7168,	2048,	 384,	5888,	-5312,	7552,	4736,	
-4032,	-5504,	-6592,	-4736,	8896,	3840,	-5824,	2240,	
-1472,	-192,	-320,	 896,	1728,	-4608,	-1856,	4288,	
1024,	-1792,	4992,	-7552,	-2752,	-6464,	-4288,	1664,	
2304,	-2368,	-4992,	-6912,	4992,	9536,	-4352,	7360,	
-4160,	-2240,	-512,	-11200,	 256,	2048,	-3264,	6912
			};

			@cb;
			@cb;
			@cb;
			@cb;
			@cb;
			go <= 1;
			@cb;
			go <= 0;
			@cb;
		
			repeat(128) @cb;
		
		for (int p=`START_POS; p>=0; p--) begin
			@cb;
			@cb;
		
			plane_start <= 1;
			bit_pos<= p;
			@cb;
			plane_start <= 0;
			@cb;
			@cb;
			for(int row = 0; row < `CB_WIDTH/4 ; row++) 
				for(int col = 0; col < `CB_WIDTH; col = col+1) begin
					first_row <= row == 0;
					second_row <= row==1;
					last_row <= row == `CB_WIDTH-1;
					one_plus_row <= row == `TILE_WIDTH/2;
					en <= 1;
					row_start <= col == 0;
					row_end <= col == `CB_WIDTH-1;
					x0 <= src[row*4  ][col][31]? (0 - src[row*4  ][col]/64) | 1<<`W_WT1 : src[row*4  ][col]/64;
					x1 <= src[row*4+1][col][31]? (0 - src[row*4+1][col]/64) | 1<<`W_WT1 : src[row*4+1][col]/64;
					x2 <= src[row*4+2][col][31]? (0 - src[row*4+2][col]/64) | 1<<`W_WT1 : src[row*4+2][col]/64;
					x3 <= src[row*4+3][col][31]? (0 - src[row*4+3][col]/64) | 1<<`W_WT1 : src[row*4+3][col]/64;
					
					@cb;
				end
			first_row <= 0;
			second_row <= 0;		
			last_row <= 0;
			one_plus_row <= 0;
			row_start <= 0;
			row_end <= 0;
			en <= 0;
			@cb;
			@cb;
			@cb;
			@cb;
			@cb;
			plane_end <= 1;
			@cb;
			plane_end <= 0;
			@cb;
			@cb;
			@cb;
			@mq_ready;
			@cb;
			repeat(11) @cb;

		end
	endtask
	
endinterface
